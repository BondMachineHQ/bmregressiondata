
`timescale 1ns/1ps
module a0(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [7:0] rom_value;


	p0 p0_instance(clock_signal, reset_signal, rom_bus, rom_value, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p0rom p0rom_instance(rom_bus, rom_value);

endmodule
`timescale 1ns/1ps
module a10(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a10din;
	wire [31:0] a10dout;
	wire [1:0] a10addr;
	wire a10wren;
	wire a10en;

	p10 p10_instance(clock_signal, reset_signal, rom_bus, rom_value, a10din, a10dout, a10addr, a10wren, a10en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p10rom p10rom_instance(rom_bus, rom_value);
	p10ram p10ram_instance(clock_signal, reset_signal, a10din, a10dout, a10addr, a10wren, a10en);

endmodule
`timescale 1ns/1ps
module a11(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a11din;
	wire [31:0] a11dout;
	wire [1:0] a11addr;
	wire a11wren;
	wire a11en;

	p11 p11_instance(clock_signal, reset_signal, rom_bus, rom_value, a11din, a11dout, a11addr, a11wren, a11en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p11rom p11rom_instance(rom_bus, rom_value);
	p11ram p11ram_instance(clock_signal, reset_signal, a11din, a11dout, a11addr, a11wren, a11en);

endmodule
`timescale 1ns/1ps
module a12(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a12din;
	wire [31:0] a12dout;
	wire [1:0] a12addr;
	wire a12wren;
	wire a12en;

	p12 p12_instance(clock_signal, reset_signal, rom_bus, rom_value, a12din, a12dout, a12addr, a12wren, a12en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p12rom p12rom_instance(rom_bus, rom_value);
	p12ram p12ram_instance(clock_signal, reset_signal, a12din, a12dout, a12addr, a12wren, a12en);

endmodule
`timescale 1ns/1ps
module a13(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a13din;
	wire [31:0] a13dout;
	wire [1:0] a13addr;
	wire a13wren;
	wire a13en;

	p13 p13_instance(clock_signal, reset_signal, rom_bus, rom_value, a13din, a13dout, a13addr, a13wren, a13en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p13rom p13rom_instance(rom_bus, rom_value);
	p13ram p13ram_instance(clock_signal, reset_signal, a13din, a13dout, a13addr, a13wren, a13en);

endmodule
`timescale 1ns/1ps
module a14(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a14din;
	wire [31:0] a14dout;
	wire [1:0] a14addr;
	wire a14wren;
	wire a14en;

	p14 p14_instance(clock_signal, reset_signal, rom_bus, rom_value, a14din, a14dout, a14addr, a14wren, a14en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p14rom p14rom_instance(rom_bus, rom_value);
	p14ram p14ram_instance(clock_signal, reset_signal, a14din, a14dout, a14addr, a14wren, a14en);

endmodule
`timescale 1ns/1ps
module a15(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a15din;
	wire [31:0] a15dout;
	wire [1:0] a15addr;
	wire a15wren;
	wire a15en;

	p15 p15_instance(clock_signal, reset_signal, rom_bus, rom_value, a15din, a15dout, a15addr, a15wren, a15en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p15rom p15rom_instance(rom_bus, rom_value);
	p15ram p15ram_instance(clock_signal, reset_signal, a15din, a15dout, a15addr, a15wren, a15en);

endmodule
`timescale 1ns/1ps
module a16(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a16din;
	wire [31:0] a16dout;
	wire [1:0] a16addr;
	wire a16wren;
	wire a16en;

	p16 p16_instance(clock_signal, reset_signal, rom_bus, rom_value, a16din, a16dout, a16addr, a16wren, a16en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p16rom p16rom_instance(rom_bus, rom_value);
	p16ram p16ram_instance(clock_signal, reset_signal, a16din, a16dout, a16addr, a16wren, a16en);

endmodule
`timescale 1ns/1ps
module a17(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a17din;
	wire [31:0] a17dout;
	wire [1:0] a17addr;
	wire a17wren;
	wire a17en;

	p17 p17_instance(clock_signal, reset_signal, rom_bus, rom_value, a17din, a17dout, a17addr, a17wren, a17en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p17rom p17rom_instance(rom_bus, rom_value);
	p17ram p17ram_instance(clock_signal, reset_signal, a17din, a17dout, a17addr, a17wren, a17en);

endmodule
`timescale 1ns/1ps
module a18(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a18din;
	wire [31:0] a18dout;
	wire [1:0] a18addr;
	wire a18wren;
	wire a18en;

	p18 p18_instance(clock_signal, reset_signal, rom_bus, rom_value, a18din, a18dout, a18addr, a18wren, a18en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p18rom p18rom_instance(rom_bus, rom_value);
	p18ram p18ram_instance(clock_signal, reset_signal, a18din, a18dout, a18addr, a18wren, a18en);

endmodule
`timescale 1ns/1ps
module a19(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a19din;
	wire [31:0] a19dout;
	wire [1:0] a19addr;
	wire a19wren;
	wire a19en;

	p19 p19_instance(clock_signal, reset_signal, rom_bus, rom_value, a19din, a19dout, a19addr, a19wren, a19en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p19rom p19rom_instance(rom_bus, rom_value);
	p19ram p19ram_instance(clock_signal, reset_signal, a19din, a19dout, a19addr, a19wren, a19en);

endmodule
`timescale 1ns/1ps
module a1(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [7:0] rom_value;


	p1 p1_instance(clock_signal, reset_signal, rom_bus, rom_value, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p1rom p1rom_instance(rom_bus, rom_value);

endmodule
`timescale 1ns/1ps
module a20(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a20din;
	wire [31:0] a20dout;
	wire [1:0] a20addr;
	wire a20wren;
	wire a20en;

	p20 p20_instance(clock_signal, reset_signal, rom_bus, rom_value, a20din, a20dout, a20addr, a20wren, a20en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p20rom p20rom_instance(rom_bus, rom_value);
	p20ram p20ram_instance(clock_signal, reset_signal, a20din, a20dout, a20addr, a20wren, a20en);

endmodule
`timescale 1ns/1ps
module a2(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [7:0] rom_value;


	p2 p2_instance(clock_signal, reset_signal, rom_bus, rom_value, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p2rom p2rom_instance(rom_bus, rom_value);

endmodule
`timescale 1ns/1ps
module a3(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [7:0] rom_value;


	p3 p3_instance(clock_signal, reset_signal, rom_bus, rom_value, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p3rom p3rom_instance(rom_bus, rom_value);

endmodule
`timescale 1ns/1ps
module a4(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, i8, i8_valid , i8_received, i9, i9_valid , i9_received, i10, i10_valid , i10_received, i11, i11_valid , i11_received, i12, i12_valid , i12_received, i13, i13_valid , i13_received, i14, i14_valid , i14_received, i15, i15_valid , i15_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received, o2, o2_valid, o2_received, o3, o3_valid, o3_received, o4, o4_valid, o4_received, o5, o5_valid, o5_received, o6, o6_valid, o6_received, o7, o7_valid, o7_received, o8, o8_valid, o8_received, o9, o9_valid, o9_received, o10, o10_valid, o10_received, o11, o11_valid, o11_received, o12, o12_valid, o12_received, o13, o13_valid, o13_received, o14, o14_valid, o14_received, o15, o15_valid, o15_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	input [31:0] i8;
	input i8_valid;
	output i8_received;
	input [31:0] i9;
	input i9_valid;
	output i9_received;
	input [31:0] i10;
	input i10_valid;
	output i10_received;
	input [31:0] i11;
	input i11_valid;
	output i11_received;
	input [31:0] i12;
	input i12_valid;
	output i12_received;
	input [31:0] i13;
	input i13_valid;
	output i13_received;
	input [31:0] i14;
	input i14_valid;
	output i14_received;
	input [31:0] i15;
	input i15_valid;
	output i15_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;
	output [31:0] o2;
	output o2_valid;
	input o2_received;
	output [31:0] o3;
	output o3_valid;
	input o3_received;
	output [31:0] o4;
	output o4_valid;
	input o4_received;
	output [31:0] o5;
	output o5_valid;
	input o5_received;
	output [31:0] o6;
	output o6_valid;
	input o6_received;
	output [31:0] o7;
	output o7_valid;
	input o7_received;
	output [31:0] o8;
	output o8_valid;
	input o8_received;
	output [31:0] o9;
	output o9_valid;
	input o9_received;
	output [31:0] o10;
	output o10_valid;
	input o10_received;
	output [31:0] o11;
	output o11_valid;
	input o11_received;
	output [31:0] o12;
	output o12_valid;
	input o12_received;
	output [31:0] o13;
	output o13_valid;
	input o13_received;
	output [31:0] o14;
	output o14_valid;
	input o14_received;
	output [31:0] o15;
	output o15_valid;
	input o15_received;

	wire [6:0] rom_bus;
	wire [37:0] rom_value;

	wire [31:0] a4din;
	wire [31:0] a4dout;
	wire [2:0] a4addr;
	wire a4wren;
	wire a4en;

	p4 p4_instance(clock_signal, reset_signal, rom_bus, rom_value, a4din, a4dout, a4addr, a4wren, a4en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, i2, i2_valid , i2_received, i3, i3_valid , i3_received, i4, i4_valid , i4_received, i5, i5_valid , i5_received, i6, i6_valid , i6_received, i7, i7_valid , i7_received, i8, i8_valid , i8_received, i9, i9_valid , i9_received, i10, i10_valid , i10_received, i11, i11_valid , i11_received, i12, i12_valid , i12_received, i13, i13_valid , i13_received, i14, i14_valid , i14_received, i15, i15_valid , i15_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received, o2, o2_valid, o2_received, o3, o3_valid, o3_received, o4, o4_valid, o4_received, o5, o5_valid, o5_received, o6, o6_valid, o6_received, o7, o7_valid, o7_received, o8, o8_valid, o8_received, o9, o9_valid, o9_received, o10, o10_valid, o10_received, o11, o11_valid, o11_received, o12, o12_valid, o12_received, o13, o13_valid, o13_received, o14, o14_valid, o14_received, o15, o15_valid, o15_received);
	p4rom p4rom_instance(rom_bus, rom_value);
	p4ram p4ram_instance(clock_signal, reset_signal, a4din, a4dout, a4addr, a4wren, a4en);

endmodule
`timescale 1ns/1ps
module a5(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a5din;
	wire [31:0] a5dout;
	wire [1:0] a5addr;
	wire a5wren;
	wire a5en;

	p5 p5_instance(clock_signal, reset_signal, rom_bus, rom_value, a5din, a5dout, a5addr, a5wren, a5en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p5rom p5rom_instance(rom_bus, rom_value);
	p5ram p5ram_instance(clock_signal, reset_signal, a5din, a5dout, a5addr, a5wren, a5en);

endmodule
`timescale 1ns/1ps
module a6(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a6din;
	wire [31:0] a6dout;
	wire [1:0] a6addr;
	wire a6wren;
	wire a6en;

	p6 p6_instance(clock_signal, reset_signal, rom_bus, rom_value, a6din, a6dout, a6addr, a6wren, a6en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p6rom p6rom_instance(rom_bus, rom_value);
	p6ram p6ram_instance(clock_signal, reset_signal, a6din, a6dout, a6addr, a6wren, a6en);

endmodule
`timescale 1ns/1ps
module a7(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a7din;
	wire [31:0] a7dout;
	wire [1:0] a7addr;
	wire a7wren;
	wire a7en;

	p7 p7_instance(clock_signal, reset_signal, rom_bus, rom_value, a7din, a7dout, a7addr, a7wren, a7en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p7rom p7rom_instance(rom_bus, rom_value);
	p7ram p7ram_instance(clock_signal, reset_signal, a7din, a7dout, a7addr, a7wren, a7en);

endmodule
`timescale 1ns/1ps
module a8(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a8din;
	wire [31:0] a8dout;
	wire [1:0] a8addr;
	wire a8wren;
	wire a8en;

	p8 p8_instance(clock_signal, reset_signal, rom_bus, rom_value, a8din, a8dout, a8addr, a8wren, a8en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p8rom p8rom_instance(rom_bus, rom_value);
	p8ram p8ram_instance(clock_signal, reset_signal, a8din, a8dout, a8addr, a8wren, a8en);

endmodule
`timescale 1ns/1ps
module a9(clock_signal, reset_signal, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

	wire [4:0] rom_bus;
	wire [38:0] rom_value;

	wire [31:0] a9din;
	wire [31:0] a9dout;
	wire [1:0] a9addr;
	wire a9wren;
	wire a9en;

	p9 p9_instance(clock_signal, reset_signal, rom_bus, rom_value, a9din, a9dout, a9addr, a9wren, a9en, i0, i0_valid , i0_received, i1, i1_valid , i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);
	p9rom p9rom_instance(rom_bus, rom_value);
	p9ram p9ram_instance(clock_signal, reset_signal, a9din, a9dout, a9addr, a9wren, a9en);

endmodule


	module bmaccelerator_v1_0 #
	(
		parameter integer C_S00_AXIS_TDATA_WIDTH	= 32,
		parameter integer C_M00_AXIS_TDATA_WIDTH	= 32,
		parameter integer C_M00_AXIS_START_COUNT	= 32
	)
	(

		input wire  s00_axis_aclk,
		input wire  s00_axis_aresetn,
		output wire  s00_axis_tready,
		input wire [C_S00_AXIS_TDATA_WIDTH-1 : 0] s00_axis_tdata,
		input wire  s00_axis_tlast,
		input wire  s00_axis_tvalid,

		input wire  m00_axis_aclk,
		input wire  m00_axis_aresetn,
		output wire  m00_axis_tvalid,
		output wire [C_M00_AXIS_TDATA_WIDTH-1 : 0] m00_axis_tdata,
		output wire  m00_axis_tlast,
		input wire  m00_axis_tready
	);


    /*
        NOW START THE AXIS SLAVE SECTION
    */

    localparam samples = 16; // number of samples that I expect from the client
    localparam bminputs = 8;  // number of bminputs for each sample (or bminputs)
    localparam bmoutputs = 8; // number of output for the classification
	localparam NUMBER_OF_INPUTS  = samples*bminputs;                                     
    localparam NUMBER_OF_OUTPUTS = samples*bmoutputs;
	localparam precision = 32; // precision bit
	localparam maxfifoloop = (C_S00_AXIS_TDATA_WIDTH / precision) - 1;
    
	// Machine state for the slave stream part
	parameter [1:0] IDLE = 1'b0,
	                WRITE_FIFO  = 1'b1; 

	wire  	   axis_tready;
	reg        mst_exec_state;     
	wire       fifo_wren;
	reg        fifo_full_flag;
	reg [11:0] write_pointer;
	reg        writes_done;
    wire       test;

	assign s00_axis_tready	= axis_tready;

	always @(posedge s00_axis_aclk) 
	begin  
	  if (!s00_axis_aresetn) 
	    begin
	      mst_exec_state <= IDLE;
	    end  
	  else
	    case (mst_exec_state)
	      IDLE:
	          if (s00_axis_tvalid)
	            begin
	              mst_exec_state <= WRITE_FIFO;
	            end
	          else
	            begin
	              mst_exec_state <= IDLE;
	            end
	      WRITE_FIFO:
	        if (writes_done)
	          begin
	            mst_exec_state <= IDLE;
	          end
	        else
	          begin
	            mst_exec_state <= WRITE_FIFO;
	          end

	    endcase
	end

	assign axis_tready = ((mst_exec_state == WRITE_FIFO) && (write_pointer <= (NUMBER_OF_INPUTS/(maxfifoloop+1))-1));

	always@(posedge s00_axis_aclk)
	begin

	  if (tx_done) begin
	       write_pointer <= 0;
	       writes_done <= 1'b0;
	  end
	  else begin
	  if(!s00_axis_aresetn)
	    begin
	      write_pointer <= 0;
	      writes_done <= 1'b0;
	    end  
	  else
	    if (write_pointer <= (NUMBER_OF_INPUTS/(maxfifoloop+1))-1)
	      begin
	        if (fifo_wren)
	          begin
	            write_pointer <= write_pointer + 1;
	            writes_done <= 1'b0;
	          end
	          if ((write_pointer == (NUMBER_OF_INPUTS/(maxfifoloop+1))-1)|| s00_axis_tlast)
	            begin
	              writes_done <= 1'b1;
	            end
	      end
	      end
	end 


	assign fifo_wren = s00_axis_tvalid && axis_tready;

	reg  [11:0] maxfifoloopcounter = 0;
	reg  [(precision)-1:0] stream_data_fifo [0 : NUMBER_OF_INPUTS-1];

	reg  [(C_S00_AXIS_TDATA_WIDTH)-1:0] stream_data_fifo [0 : NUMBER_OF_INPUTS-1];
    always @( posedge s00_axis_aclk )
    begin
		if (tx_done) begin
	       maxfifoloopcounter <= 0;
	  end
      if (fifo_wren)
        begin
          if (precision == 32) begin
            stream_data_fifo[write_pointer+maxfifoloopcounter] <= s00_axis_tdata;
            maxfifoloopcounter <= maxfifoloopcounter + 0;
          end
          else if (precision == 16) begin
              stream_data_fifo[write_pointer+maxfifoloopcounter+0] <= s00_axis_tdata[15:0];
              stream_data_fifo[write_pointer+maxfifoloopcounter+1] <= s00_axis_tdata[31:16];
              maxfifoloopcounter <= maxfifoloopcounter + 1;
          end
        end   
     end      

    /*
        NOW START THE MASTER AXIS SECTION
    */
                             
	parameter [1:0] IDLE_M = 2'b00,                                             
	                INIT_COUNTER_M  = 2'b01, 
	                PROCESS_BM = 2'B10,   
	                SEND_STREAM_M   = 2'b11; 

	reg [1:0]   mst_exec_state_M;
    reg [11:0] 	count;

    wire  	axis_tvalid;
    reg  	axis_tvalid_delay;
    wire  	axis_tlast;
    reg  	axis_tlast_delay;
    reg [C_M00_AXIS_TDATA_WIDTH-1 : 0] 	stream_data_out;
    wire  	tx_en;
    reg  	tx_done;
    wire     bm_done;

    reg  [11:0] outputs_counter = 0;
    reg  [11:0] outputs_counter_incr = 0;
	reg  [11:0] outputs_counter_pointer = 0;
    reg  [11:0] stream_output_counter = 0;
    reg  [(C_S00_AXIS_TDATA_WIDTH)-1:0] output_stream_data_fifo [0 : NUMBER_OF_OUTPUTS-1];

    assign m00_axis_tvalid	= axis_tvalid_delay;
	assign m00_axis_tdata	= stream_data_out;
	assign m00_axis_tlast	= axis_tlast_delay;

	always @(posedge m00_axis_aclk)                                             
	begin                                                                     
	  if (!m00_axis_aresetn)                                                  
	    begin                                                                 
	      mst_exec_state_M <= IDLE_M;                                             
	      count    <= 0;                                                      
	    end                                                                   
	  else                                                                    
	    case (mst_exec_state_M)                                                 
	      IDLE_M:                                                         
	            mst_exec_state_M  <= INIT_COUNTER_M; 

	      INIT_COUNTER_M:                              
	        if ( count == 32 - 1 )                               
	          begin                                                           
	            mst_exec_state_M  <= PROCESS_BM;                               
	          end                                                             
	        else                                                              
	          begin                                                           
	            count <= count + 1;                                           
	            mst_exec_state_M  <= INIT_COUNTER_M;                              
	          end                                                             

	      PROCESS_BM:
	           if (!bm_done) 
	           begin
	               mst_exec_state_M <= PROCESS_BM;
	           end
	           else
	           begin
	               mst_exec_state_M <= SEND_STREAM_M;   
	           end

	      SEND_STREAM_M:                          
	        if (tx_done)                                                      
	          begin                                                           
	            mst_exec_state_M <= IDLE_M;                                       
	          end                                                             
	        else                                                              
	          begin                                                           
	            mst_exec_state_M <= SEND_STREAM_M;                                
	          end                                                             
	    endcase                                                               
	end

	assign axis_tvalid = ((mst_exec_state_M == SEND_STREAM_M) && (writes_done) && (bm_done));
    assign axis_tlast = (stream_output_counter == (NUMBER_OF_OUTPUTS/(maxfifoloop+1)) - 1);

    always @(posedge m00_axis_aclk)                                                                  
	begin        
	if (tx_done) begin
	       axis_tvalid_delay <= 1'b0;                                                               
	      axis_tlast_delay <= 1'b0;         
	end     
	else begin                                                                             
	  if (!m00_axis_aresetn)                                                                         
	    begin                                                                                      
	      axis_tvalid_delay <= 1'b0;                                                               
	      axis_tlast_delay <= 1'b0;                                                                
	    end                                                                                        
	  else                                                                                         
	    begin                                                                                      
	      axis_tvalid_delay <= axis_tvalid;                                                        
	      axis_tlast_delay <= axis_tlast;                                                          
	    end                                                                                        
	end 
	end
	reg [31:0] i0_r = 32'b0;
	reg [31:0] i1_r = 32'b0;
	reg [31:0] i2_r = 32'b0;
	reg [31:0] i3_r = 32'b0;
	reg [31:0] i4_r = 32'b0;
	reg [31:0] i5_r = 32'b0;
	reg [31:0] i6_r = 32'b0;
	reg [31:0] i7_r = 32'b0;
	reg [31:0] o0_received_r;
	reg [31:0] o1_received_r;
	reg [31:0] o2_received_r;
	reg [31:0] o3_received_r;
	reg [31:0] o4_received_r;
	reg [31:0] o5_received_r;
	reg [31:0] o6_received_r;
	reg [31:0] o7_received_r;
	wire [31:0] i0;
	wire i0_valid;
	wire i0_received;
	wire [31:0] i1;
	wire i1_valid;
	wire i1_received;
	wire [31:0] i2;
	wire i2_valid;
	wire i2_received;
	wire [31:0] i3;
	wire i3_valid;
	wire i3_received;
	wire [31:0] i4;
	wire i4_valid;
	wire i4_received;
	wire [31:0] i5;
	wire i5_valid;
	wire i5_received;
	wire [31:0] i6;
	wire i6_valid;
	wire i6_received;
	wire [31:0] i7;
	wire i7_valid;
	wire i7_received;
	reg i0_valid_r = 1'b0;
	reg i1_valid_r = 1'b0;
	reg i2_valid_r = 1'b0;
	reg i3_valid_r = 1'b0;
	reg i4_valid_r = 1'b0;
	reg i5_valid_r = 1'b0;
	reg i6_valid_r = 1'b0;
	reg i7_valid_r = 1'b0;
	wire [31:0] o0;
	wire o0_valid;
	wire o0_received;
	reg  o0_valid_r = 1'b0;
	wire [31:0] o1;
	wire o1_valid;
	wire o1_received;
	reg  o1_valid_r = 1'b0;
	wire [31:0] o2;
	wire o2_valid;
	wire o2_received;
	reg  o2_valid_r = 1'b0;
	wire [31:0] o3;
	wire o3_valid;
	wire o3_received;
	reg  o3_valid_r = 1'b0;
	wire [31:0] o4;
	wire o4_valid;
	wire o4_received;
	reg  o4_valid_r = 1'b0;
	wire [31:0] o5;
	wire o5_valid;
	wire o5_received;
	reg  o5_valid_r = 1'b0;
	wire [31:0] o6;
	wire o6_valid;
	wire o6_received;
	reg  o6_valid_r = 1'b0;
	wire [31:0] o7;
	wire o7_valid;
	wire o7_received;
	reg  o7_valid_r = 1'b0;
	assign i0 = i0_r;
	assign i1 = i1_r;
	assign i2 = i2_r;
	assign i3 = i3_r;
	assign i4 = i4_r;
	assign i5 = i5_r;
	assign i6 = i6_r;
	assign i7 = i7_r;
	assign i0_valid = i0_valid_r;
	assign i1_valid = i1_valid_r;
	assign i2_valid = i2_valid_r;
	assign i3_valid = i3_valid_r;
	assign i4_valid = i4_valid_r;
	assign i5_valid = i5_valid_r;
	assign i6_valid = i6_valid_r;
	assign i7_valid = i7_valid_r;
	assign o0_received = o0_received_r;
	assign o1_received = o1_received_r;
	assign o2_received = o2_received_r;
	assign o3_received = o3_received_r;
	assign o4_received = o4_received_r;
	assign o5_received = o5_received_r;
	assign o6_received = o6_received_r;
	assign o7_received = o7_received_r;

    assign bm_done = (outputs_counter_incr == samples);
	reg[1:0] send = 2'b00;

	bondmachine bm(.clk(m00_axis_aclk),
	.reset(!m00_axis_aresetn),
	.i0(i0),
	.i0_valid(i0_valid),
	.i0_received(i0_received),
	.i1(i1),
	.i1_valid(i1_valid),
	.i1_received(i1_received),
	.i2(i2),
	.i2_valid(i2_valid),
	.i2_received(i2_received),
	.i3(i3),
	.i3_valid(i3_valid),
	.i3_received(i3_received),
	.i4(i4),
	.i4_valid(i4_valid),
	.i4_received(i4_received),
	.i5(i5),
	.i5_valid(i5_valid),
	.i5_received(i5_received),
	.i6(i6),
	.i6_valid(i6_valid),
	.i6_received(i6_received),
	.i7(i7),
	.i7_valid(i7_valid),
	.i7_received(i7_received),
	.o0(o0),
	.o0_valid(o0_valid),
	.o0_received(o0_received),
	.o1(o1),
	.o1_valid(o1_valid),
	.o1_received(o1_received),
	.o2(o2),
	.o2_valid(o2_valid),
	.o2_received(o2_received),
	.o3(o3),
	.o3_valid(o3_valid),
	.o3_received(o3_received),
	.o4(o4),
	.o4_valid(o4_valid),
	.o4_received(o4_received),
	.o5(o5),
	.o5_valid(o5_valid),
	.o5_received(o5_received),
	.o6(o6),
	.o6_valid(o6_valid),
	.o6_received(o6_received),
	.o7(o7),
	.o7_valid(o7_valid),
	.o7_received(o7_received)
	);

    always @( posedge m00_axis_aclk )                  
	begin        
    
        if (tx_done) begin
            outputs_counter <= 0;
            outputs_counter_incr <= 0;
			outputs_counter_pointer <= 0;
			o0_received_r <= 1'b0;
			o0_valid_r <= 1'b0;
			o1_received_r <= 1'b0;
			o1_valid_r <= 1'b0;
			o2_received_r <= 1'b0;
			o2_valid_r <= 1'b0;
			o3_received_r <= 1'b0;
			o3_valid_r <= 1'b0;
			o4_received_r <= 1'b0;
			o4_valid_r <= 1'b0;
			o5_received_r <= 1'b0;
			o5_valid_r <= 1'b0;
			o6_received_r <= 1'b0;
			o6_valid_r <= 1'b0;
			o7_received_r <= 1'b0;
			o7_valid_r <= 1'b0;
        end
        else begin
            if (writes_done && !bm_done) begin
            
			if (send == 2'b00) begin
				send <= 2'b01;
				i0_r <= stream_data_fifo[outputs_counter+0];
				i1_r <= stream_data_fifo[outputs_counter+1];
				i2_r <= stream_data_fifo[outputs_counter+2];
				i3_r <= stream_data_fifo[outputs_counter+3];
				i4_r <= stream_data_fifo[outputs_counter+4];
				i5_r <= stream_data_fifo[outputs_counter+5];
				i6_r <= stream_data_fifo[outputs_counter+6];
				i7_r <= stream_data_fifo[outputs_counter+7];
				i0_valid_r <= 1'b1;
				i1_valid_r <= 1'b1;
				i2_valid_r <= 1'b1;
				i3_valid_r <= 1'b1;
				i4_valid_r <= 1'b1;
				i5_valid_r <= 1'b1;
				i6_valid_r <= 1'b1;
				i7_valid_r <= 1'b1;
			end
			else if (send == 2'b01) begin
			    if (
					i0_received &&
					i1_received &&
					i2_received &&
					i3_received &&
					i4_received &&
					i5_received &&
					i6_received &&
					i7_received
				) begin
					i0_valid_r <= 1'b0;
					i1_valid_r <= 1'b0;
					i2_valid_r <= 1'b0;
					i3_valid_r <= 1'b0;
					i4_valid_r <= 1'b0;
					i5_valid_r <= 1'b0;
					i6_valid_r <= 1'b0;
					i7_valid_r <= 1'b0;

					send <= 2'b10;
				end
			end
			else if (send == 2'b10) begin
			if ( o0_valid && !o0_received_r) begin
				o0_valid_r <= 1'b1;
				o0_received_r <= 1'b1;
				output_stream_data_fifo[outputs_counter_pointer+0] <= o0;
			end
			if ( o1_valid && !o1_received_r) begin
				o1_valid_r <= 1'b1;
				o1_received_r <= 1'b1;
				output_stream_data_fifo[outputs_counter_pointer+1] <= o1;
			end
			if ( o2_valid && !o2_received_r) begin
				o2_valid_r <= 1'b1;
				o2_received_r <= 1'b1;
				output_stream_data_fifo[outputs_counter_pointer+2] <= o2;
			end
			if ( o3_valid && !o3_received_r) begin
				o3_valid_r <= 1'b1;
				o3_received_r <= 1'b1;
				output_stream_data_fifo[outputs_counter_pointer+3] <= o3;
			end
			if ( o4_valid && !o4_received_r) begin
				o4_valid_r <= 1'b1;
				o4_received_r <= 1'b1;
				output_stream_data_fifo[outputs_counter_pointer+4] <= o4;
			end
			if ( o5_valid && !o5_received_r) begin
				o5_valid_r <= 1'b1;
				o5_received_r <= 1'b1;
				output_stream_data_fifo[outputs_counter_pointer+5] <= o5;
			end
			if ( o6_valid && !o6_received_r) begin
				o6_valid_r <= 1'b1;
				o6_received_r <= 1'b1;
				output_stream_data_fifo[outputs_counter_pointer+6] <= o6;
			end
			if ( o7_valid && !o7_received_r) begin
				o7_valid_r <= 1'b1;
				o7_received_r <= 1'b1;
				output_stream_data_fifo[outputs_counter_pointer+7] <= o7;
			end

			if (
				o0_valid_r &&
				o1_valid_r &&
				o2_valid_r &&
				o3_valid_r &&
				o4_valid_r &&
				o5_valid_r &&
				o6_valid_r &&
				o7_valid_r

			 ) begin
				o0_valid_r <= 1'b0;
				o1_valid_r <= 1'b0;
				o2_valid_r <= 1'b0;
				o3_valid_r <= 1'b0;
				o4_valid_r <= 1'b0;
				o5_valid_r <= 1'b0;
				o6_valid_r <= 1'b0;
				o7_valid_r <= 1'b0;

			end
			else if(
				!o0_valid && o0_received_r &&
				!o1_valid && o1_received_r &&
				!o2_valid && o2_received_r &&
				!o3_valid && o3_received_r &&
				!o4_valid && o4_received_r &&
				!o5_valid && o5_received_r &&
				!o6_valid && o6_received_r &&
				!o7_valid && o7_received_r
			) 
			begin
					o0_received_r <= 1'b0;
					o1_received_r <= 1'b0;
					o2_received_r <= 1'b0;
					o3_received_r <= 1'b0;
					o4_received_r <= 1'b0;
					o5_received_r <= 1'b0;
					o6_received_r <= 1'b0;
					o7_received_r <= 1'b0;
					outputs_counter_pointer <= outputs_counter_pointer + bmoutputs;
					outputs_counter_incr <= outputs_counter_incr + 1;
					outputs_counter <= bminputs*(outputs_counter_incr+1);
					
					send <= 2'b00;
			end
			end
			end
	    end
	end

    assign tx_en = m00_axis_tready && axis_tvalid;   

	reg [11:0] maxfifoloopcounteroutput = 0;

    always @( posedge m00_axis_aclk )                  
    begin        
       if (tx_done) begin
		maxfifoloopcounteroutput <= 0;
        stream_output_counter <= 0;
        tx_done <= 1'b0;
       end
                                     
      if(!m00_axis_aresetn)                            
        begin   
          stream_data_out <= 1;                      
        end                                          
      else if (tx_en)
        begin
           if (stream_output_counter <= (NUMBER_OF_OUTPUTS/(maxfifoloop+1)) - 1) begin
              if (precision == 32) begin
                    stream_data_out <= output_stream_data_fifo[stream_output_counter+maxfifoloopcounteroutput];
              end
              else if (precision == 16) begin
                    //stream_data_out <= output_stream_data_fifo[stream_output_counter+maxfifoloopcounteroutput];
                    stream_data_out[15:0] <= output_stream_data_fifo[stream_output_counter+maxfifoloopcounteroutput+0];
                    stream_data_out[31:16] <= output_stream_data_fifo[stream_output_counter+maxfifoloopcounteroutput+1];
                    maxfifoloopcounteroutput <= maxfifoloopcounteroutput + 1;
              end
              stream_output_counter <= stream_output_counter + 1;
              if (stream_output_counter == (NUMBER_OF_OUTPUTS/(maxfifoloop+1)) - 1) begin
                    tx_done <= 1'b1;
              end
          end
        end                                          
    end

endmodule

module bondmachine(clk, reset, i0, i0_valid, i0_received, i1, i1_valid, i1_received, i2, i2_valid, i2_received, i3, i3_valid, i3_received, i4, i4_valid, i4_received, i5, i5_valid, i5_received, i6, i6_valid, i6_received, i7, i7_valid, i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received, o2, o2_valid, o2_received, o3, o3_valid, o3_received, o4, o4_valid, o4_received, o5, o5_valid, o5_received, o6, o6_valid, o6_received, o7, o7_valid, o7_received);

	// Clock and reset input ports
	input clk, reset;
	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	//--------------Output Ports-----------------------
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;
	output [31:0] o2;
	output o2_valid;
	input o2_received;
	output [31:0] o3;
	output o3_valid;
	input o3_received;
	output [31:0] o4;
	output o4_valid;
	input o4_received;
	output [31:0] o5;
	output o5_valid;
	input o5_received;
	output [31:0] o6;
	output o6_valid;
	input o6_received;
	output [31:0] o7;
	output o7_valid;
	input o7_received;



	//Analyzing Internal output p0o0
	//Internal output p0o0 is connected to p4i8
	wire [31:0] p0o0;
	wire p0o0_valid;
	wire p0o0_received;
	wire p4i8_received;
	//Analyzing Internal output p0o1
	//Internal output p0o1 is connected to p4i9
	wire [31:0] p0o1;
	wire p0o1_valid;
	wire p0o1_received;
	wire p4i9_received;
	//Analyzing Internal output p1o0
	//Internal output p1o0 is connected to p4i10
	wire [31:0] p1o0;
	wire p1o0_valid;
	wire p1o0_received;
	wire p4i10_received;
	//Analyzing Internal output p1o1
	//Internal output p1o1 is connected to p4i11
	wire [31:0] p1o1;
	wire p1o1_valid;
	wire p1o1_received;
	wire p4i11_received;
	//Analyzing Internal output p2o0
	//Internal output p2o0 is connected to p4i12
	wire [31:0] p2o0;
	wire p2o0_valid;
	wire p2o0_received;
	wire p4i12_received;
	//Analyzing Internal output p2o1
	//Internal output p2o1 is connected to p4i13
	wire [31:0] p2o1;
	wire p2o1_valid;
	wire p2o1_received;
	wire p4i13_received;
	//Analyzing Internal output p3o0
	//Internal output p3o0 is connected to p4i14
	wire [31:0] p3o0;
	wire p3o0_valid;
	wire p3o0_received;
	wire p4i14_received;
	//Analyzing Internal output p3o1
	//Internal output p3o1 is connected to p4i15
	wire [31:0] p3o1;
	wire p3o1_valid;
	wire p3o1_received;
	wire p4i15_received;
	//Analyzing Internal output p4o0
	//Internal output p4o0 is connected to o0
	wire [31:0] p4o0;
	wire p4o0_valid;
	wire p4o0_received;
	wire o0_received;
	//Analyzing Internal output p4o1
	//Internal output p4o1 is connected to o1
	wire [31:0] p4o1;
	wire p4o1_valid;
	wire p4o1_received;
	wire o1_received;
	//Analyzing Internal output p4o2
	//Internal output p4o2 is connected to o2
	wire [31:0] p4o2;
	wire p4o2_valid;
	wire p4o2_received;
	wire o2_received;
	//Analyzing Internal output p4o3
	//Internal output p4o3 is connected to o3
	wire [31:0] p4o3;
	wire p4o3_valid;
	wire p4o3_received;
	wire o3_received;
	//Analyzing Internal output p4o4
	//Internal output p4o4 is connected to o4
	wire [31:0] p4o4;
	wire p4o4_valid;
	wire p4o4_received;
	wire o4_received;
	//Analyzing Internal output p4o5
	//Internal output p4o5 is connected to o5
	wire [31:0] p4o5;
	wire p4o5_valid;
	wire p4o5_received;
	wire o5_received;
	//Analyzing Internal output p4o6
	//Internal output p4o6 is connected to o6
	wire [31:0] p4o6;
	wire p4o6_valid;
	wire p4o6_received;
	wire o6_received;
	//Analyzing Internal output p4o7
	//Internal output p4o7 is connected to o7
	wire [31:0] p4o7;
	wire p4o7_valid;
	wire p4o7_received;
	wire o7_received;
	//Analyzing Internal output p4o8
	//Internal output p4o8 is connected to p5i0
	//Internal output p4o8 is connected to p9i0
	//Internal output p4o8 is connected to p13i0
	//Internal output p4o8 is connected to p17i0
	wire [31:0] p4o8;
	wire p4o8_valid;
	wire p4o8_received;
	wire p5i0_received;
	wire p9i0_received;
	wire p13i0_received;
	wire p17i0_received;
	//Analyzing Internal output p4o9
	//Internal output p4o9 is connected to p5i1
	//Internal output p4o9 is connected to p9i1
	//Internal output p4o9 is connected to p13i1
	//Internal output p4o9 is connected to p17i1
	wire [31:0] p4o9;
	wire p4o9_valid;
	wire p4o9_received;
	wire p5i1_received;
	wire p9i1_received;
	wire p13i1_received;
	wire p17i1_received;
	//Analyzing Internal output p4o10
	//Internal output p4o10 is connected to p6i0
	//Internal output p4o10 is connected to p10i0
	//Internal output p4o10 is connected to p14i0
	//Internal output p4o10 is connected to p18i0
	wire [31:0] p4o10;
	wire p4o10_valid;
	wire p4o10_received;
	wire p6i0_received;
	wire p10i0_received;
	wire p14i0_received;
	wire p18i0_received;
	//Analyzing Internal output p4o11
	//Internal output p4o11 is connected to p6i1
	//Internal output p4o11 is connected to p10i1
	//Internal output p4o11 is connected to p14i1
	//Internal output p4o11 is connected to p18i1
	wire [31:0] p4o11;
	wire p4o11_valid;
	wire p4o11_received;
	wire p6i1_received;
	wire p10i1_received;
	wire p14i1_received;
	wire p18i1_received;
	//Analyzing Internal output p4o12
	//Internal output p4o12 is connected to p7i0
	//Internal output p4o12 is connected to p11i0
	//Internal output p4o12 is connected to p15i0
	//Internal output p4o12 is connected to p19i0
	wire [31:0] p4o12;
	wire p4o12_valid;
	wire p4o12_received;
	wire p7i0_received;
	wire p11i0_received;
	wire p15i0_received;
	wire p19i0_received;
	//Analyzing Internal output p4o13
	//Internal output p4o13 is connected to p7i1
	//Internal output p4o13 is connected to p11i1
	//Internal output p4o13 is connected to p15i1
	//Internal output p4o13 is connected to p19i1
	wire [31:0] p4o13;
	wire p4o13_valid;
	wire p4o13_received;
	wire p7i1_received;
	wire p11i1_received;
	wire p15i1_received;
	wire p19i1_received;
	//Analyzing Internal output p4o14
	//Internal output p4o14 is connected to p8i0
	//Internal output p4o14 is connected to p12i0
	//Internal output p4o14 is connected to p16i0
	//Internal output p4o14 is connected to p20i0
	wire [31:0] p4o14;
	wire p4o14_valid;
	wire p4o14_received;
	wire p8i0_received;
	wire p12i0_received;
	wire p16i0_received;
	wire p20i0_received;
	//Analyzing Internal output p4o15
	//Internal output p4o15 is connected to p8i1
	//Internal output p4o15 is connected to p12i1
	//Internal output p4o15 is connected to p16i1
	//Internal output p4o15 is connected to p20i1
	wire [31:0] p4o15;
	wire p4o15_valid;
	wire p4o15_received;
	wire p8i1_received;
	wire p12i1_received;
	wire p16i1_received;
	wire p20i1_received;
	//Analyzing Internal output p5o0
	//Internal output p5o0 is connected to p0i0
	wire [31:0] p5o0;
	wire p5o0_valid;
	wire p5o0_received;
	wire p0i0_received;
	//Analyzing Internal output p5o1
	//Internal output p5o1 is connected to p0i1
	wire [31:0] p5o1;
	wire p5o1_valid;
	wire p5o1_received;
	wire p0i1_received;
	//Analyzing Internal output p6o0
	//Internal output p6o0 is connected to p0i2
	wire [31:0] p6o0;
	wire p6o0_valid;
	wire p6o0_received;
	wire p0i2_received;
	//Analyzing Internal output p6o1
	//Internal output p6o1 is connected to p0i3
	wire [31:0] p6o1;
	wire p6o1_valid;
	wire p6o1_received;
	wire p0i3_received;
	//Analyzing Internal output p7o0
	//Internal output p7o0 is connected to p0i4
	wire [31:0] p7o0;
	wire p7o0_valid;
	wire p7o0_received;
	wire p0i4_received;
	//Analyzing Internal output p7o1
	//Internal output p7o1 is connected to p0i5
	wire [31:0] p7o1;
	wire p7o1_valid;
	wire p7o1_received;
	wire p0i5_received;
	//Analyzing Internal output p8o0
	//Internal output p8o0 is connected to p0i6
	wire [31:0] p8o0;
	wire p8o0_valid;
	wire p8o0_received;
	wire p0i6_received;
	//Analyzing Internal output p8o1
	//Internal output p8o1 is connected to p0i7
	wire [31:0] p8o1;
	wire p8o1_valid;
	wire p8o1_received;
	wire p0i7_received;
	//Analyzing Internal output p9o0
	//Internal output p9o0 is connected to p1i0
	wire [31:0] p9o0;
	wire p9o0_valid;
	wire p9o0_received;
	wire p1i0_received;
	//Analyzing Internal output p9o1
	//Internal output p9o1 is connected to p1i1
	wire [31:0] p9o1;
	wire p9o1_valid;
	wire p9o1_received;
	wire p1i1_received;
	//Analyzing Internal output p10o0
	//Internal output p10o0 is connected to p1i2
	wire [31:0] p10o0;
	wire p10o0_valid;
	wire p10o0_received;
	wire p1i2_received;
	//Analyzing Internal output p10o1
	//Internal output p10o1 is connected to p1i3
	wire [31:0] p10o1;
	wire p10o1_valid;
	wire p10o1_received;
	wire p1i3_received;
	//Analyzing Internal output p11o0
	//Internal output p11o0 is connected to p1i4
	wire [31:0] p11o0;
	wire p11o0_valid;
	wire p11o0_received;
	wire p1i4_received;
	//Analyzing Internal output p11o1
	//Internal output p11o1 is connected to p1i5
	wire [31:0] p11o1;
	wire p11o1_valid;
	wire p11o1_received;
	wire p1i5_received;
	//Analyzing Internal output p12o0
	//Internal output p12o0 is connected to p1i6
	wire [31:0] p12o0;
	wire p12o0_valid;
	wire p12o0_received;
	wire p1i6_received;
	//Analyzing Internal output p12o1
	//Internal output p12o1 is connected to p1i7
	wire [31:0] p12o1;
	wire p12o1_valid;
	wire p12o1_received;
	wire p1i7_received;
	//Analyzing Internal output p13o0
	//Internal output p13o0 is connected to p2i0
	wire [31:0] p13o0;
	wire p13o0_valid;
	wire p13o0_received;
	wire p2i0_received;
	//Analyzing Internal output p13o1
	//Internal output p13o1 is connected to p2i1
	wire [31:0] p13o1;
	wire p13o1_valid;
	wire p13o1_received;
	wire p2i1_received;
	//Analyzing Internal output p14o0
	//Internal output p14o0 is connected to p2i2
	wire [31:0] p14o0;
	wire p14o0_valid;
	wire p14o0_received;
	wire p2i2_received;
	//Analyzing Internal output p14o1
	//Internal output p14o1 is connected to p2i3
	wire [31:0] p14o1;
	wire p14o1_valid;
	wire p14o1_received;
	wire p2i3_received;
	//Analyzing Internal output p15o0
	//Internal output p15o0 is connected to p2i4
	wire [31:0] p15o0;
	wire p15o0_valid;
	wire p15o0_received;
	wire p2i4_received;
	//Analyzing Internal output p15o1
	//Internal output p15o1 is connected to p2i5
	wire [31:0] p15o1;
	wire p15o1_valid;
	wire p15o1_received;
	wire p2i5_received;
	//Analyzing Internal output p16o0
	//Internal output p16o0 is connected to p2i6
	wire [31:0] p16o0;
	wire p16o0_valid;
	wire p16o0_received;
	wire p2i6_received;
	//Analyzing Internal output p16o1
	//Internal output p16o1 is connected to p2i7
	wire [31:0] p16o1;
	wire p16o1_valid;
	wire p16o1_received;
	wire p2i7_received;
	//Analyzing Internal output p17o0
	//Internal output p17o0 is connected to p3i0
	wire [31:0] p17o0;
	wire p17o0_valid;
	wire p17o0_received;
	wire p3i0_received;
	//Analyzing Internal output p17o1
	//Internal output p17o1 is connected to p3i1
	wire [31:0] p17o1;
	wire p17o1_valid;
	wire p17o1_received;
	wire p3i1_received;
	//Analyzing Internal output p18o0
	//Internal output p18o0 is connected to p3i2
	wire [31:0] p18o0;
	wire p18o0_valid;
	wire p18o0_received;
	wire p3i2_received;
	//Analyzing Internal output p18o1
	//Internal output p18o1 is connected to p3i3
	wire [31:0] p18o1;
	wire p18o1_valid;
	wire p18o1_received;
	wire p3i3_received;
	//Analyzing Internal output p19o0
	//Internal output p19o0 is connected to p3i4
	wire [31:0] p19o0;
	wire p19o0_valid;
	wire p19o0_received;
	wire p3i4_received;
	//Analyzing Internal output p19o1
	//Internal output p19o1 is connected to p3i5
	wire [31:0] p19o1;
	wire p19o1_valid;
	wire p19o1_received;
	wire p3i5_received;
	//Analyzing Internal output p20o0
	//Internal output p20o0 is connected to p3i6
	wire [31:0] p20o0;
	wire p20o0_valid;
	wire p20o0_received;
	wire p3i6_received;
	//Analyzing Internal output p20o1
	//Internal output p20o1 is connected to p3i7
	wire [31:0] p20o1;
	wire p20o1_valid;
	wire p20o1_received;
	wire p3i7_received;
	//Analyzing Internal output i0
	//Internal output i0 is connected to p4i0
	wire [31:0] i0;
	wire i0_valid;
	wire i0_received;
	wire p4i0_received;
	//Analyzing Internal output i1
	//Internal output i1 is connected to p4i1
	wire [31:0] i1;
	wire i1_valid;
	wire i1_received;
	wire p4i1_received;
	//Analyzing Internal output i2
	//Internal output i2 is connected to p4i2
	wire [31:0] i2;
	wire i2_valid;
	wire i2_received;
	wire p4i2_received;
	//Analyzing Internal output i3
	//Internal output i3 is connected to p4i3
	wire [31:0] i3;
	wire i3_valid;
	wire i3_received;
	wire p4i3_received;
	//Analyzing Internal output i4
	//Internal output i4 is connected to p4i4
	wire [31:0] i4;
	wire i4_valid;
	wire i4_received;
	wire p4i4_received;
	//Analyzing Internal output i5
	//Internal output i5 is connected to p4i5
	wire [31:0] i5;
	wire i5_valid;
	wire i5_received;
	wire p4i5_received;
	//Analyzing Internal output i6
	//Internal output i6 is connected to p4i6
	wire [31:0] i6;
	wire i6_valid;
	wire i6_received;
	wire p4i6_received;
	//Analyzing Internal output i7
	//Internal output i7 is connected to p4i7
	wire [31:0] i7;
	wire i7_valid;
	wire i7_received;
	wire p4i7_received;


	//Instantiation of the Processors and Shared Objects
	a0 a0_inst(clk, reset, p5o0, p5o0_valid, p0i0_received, p5o1, p5o1_valid, p0i1_received, p6o0, p6o0_valid, p0i2_received, p6o1, p6o1_valid, p0i3_received, p7o0, p7o0_valid, p0i4_received, p7o1, p7o1_valid, p0i5_received, p8o0, p8o0_valid, p0i6_received, p8o1, p8o1_valid, p0i7_received, p0o0, p0o0_valid, p0o0_received, p0o1, p0o1_valid, p0o1_received);
	a1 a1_inst(clk, reset, p9o0, p9o0_valid, p1i0_received, p9o1, p9o1_valid, p1i1_received, p10o0, p10o0_valid, p1i2_received, p10o1, p10o1_valid, p1i3_received, p11o0, p11o0_valid, p1i4_received, p11o1, p11o1_valid, p1i5_received, p12o0, p12o0_valid, p1i6_received, p12o1, p12o1_valid, p1i7_received, p1o0, p1o0_valid, p1o0_received, p1o1, p1o1_valid, p1o1_received);
	a2 a2_inst(clk, reset, p13o0, p13o0_valid, p2i0_received, p13o1, p13o1_valid, p2i1_received, p14o0, p14o0_valid, p2i2_received, p14o1, p14o1_valid, p2i3_received, p15o0, p15o0_valid, p2i4_received, p15o1, p15o1_valid, p2i5_received, p16o0, p16o0_valid, p2i6_received, p16o1, p16o1_valid, p2i7_received, p2o0, p2o0_valid, p2o0_received, p2o1, p2o1_valid, p2o1_received);
	a3 a3_inst(clk, reset, p17o0, p17o0_valid, p3i0_received, p17o1, p17o1_valid, p3i1_received, p18o0, p18o0_valid, p3i2_received, p18o1, p18o1_valid, p3i3_received, p19o0, p19o0_valid, p3i4_received, p19o1, p19o1_valid, p3i5_received, p20o0, p20o0_valid, p3i6_received, p20o1, p20o1_valid, p3i7_received, p3o0, p3o0_valid, p3o0_received, p3o1, p3o1_valid, p3o1_received);
	a4 a4_inst(clk, reset, i0, i0_valid, p4i0_received, i1, i1_valid, p4i1_received, i2, i2_valid, p4i2_received, i3, i3_valid, p4i3_received, i4, i4_valid, p4i4_received, i5, i5_valid, p4i5_received, i6, i6_valid, p4i6_received, i7, i7_valid, p4i7_received, p0o0, p0o0_valid, p4i8_received, p0o1, p0o1_valid, p4i9_received, p1o0, p1o0_valid, p4i10_received, p1o1, p1o1_valid, p4i11_received, p2o0, p2o0_valid, p4i12_received, p2o1, p2o1_valid, p4i13_received, p3o0, p3o0_valid, p4i14_received, p3o1, p3o1_valid, p4i15_received, p4o0, p4o0_valid, p4o0_received, p4o1, p4o1_valid, p4o1_received, p4o2, p4o2_valid, p4o2_received, p4o3, p4o3_valid, p4o3_received, p4o4, p4o4_valid, p4o4_received, p4o5, p4o5_valid, p4o5_received, p4o6, p4o6_valid, p4o6_received, p4o7, p4o7_valid, p4o7_received, p4o8, p4o8_valid, p4o8_received, p4o9, p4o9_valid, p4o9_received, p4o10, p4o10_valid, p4o10_received, p4o11, p4o11_valid, p4o11_received, p4o12, p4o12_valid, p4o12_received, p4o13, p4o13_valid, p4o13_received, p4o14, p4o14_valid, p4o14_received, p4o15, p4o15_valid, p4o15_received);
	a5 a5_inst(clk, reset, p4o8, p4o8_valid, p5i0_received, p4o9, p4o9_valid, p5i1_received, p5o0, p5o0_valid, p5o0_received, p5o1, p5o1_valid, p5o1_received);
	a6 a6_inst(clk, reset, p4o10, p4o10_valid, p6i0_received, p4o11, p4o11_valid, p6i1_received, p6o0, p6o0_valid, p6o0_received, p6o1, p6o1_valid, p6o1_received);
	a7 a7_inst(clk, reset, p4o12, p4o12_valid, p7i0_received, p4o13, p4o13_valid, p7i1_received, p7o0, p7o0_valid, p7o0_received, p7o1, p7o1_valid, p7o1_received);
	a8 a8_inst(clk, reset, p4o14, p4o14_valid, p8i0_received, p4o15, p4o15_valid, p8i1_received, p8o0, p8o0_valid, p8o0_received, p8o1, p8o1_valid, p8o1_received);
	a9 a9_inst(clk, reset, p4o8, p4o8_valid, p9i0_received, p4o9, p4o9_valid, p9i1_received, p9o0, p9o0_valid, p9o0_received, p9o1, p9o1_valid, p9o1_received);
	a10 a10_inst(clk, reset, p4o10, p4o10_valid, p10i0_received, p4o11, p4o11_valid, p10i1_received, p10o0, p10o0_valid, p10o0_received, p10o1, p10o1_valid, p10o1_received);
	a11 a11_inst(clk, reset, p4o12, p4o12_valid, p11i0_received, p4o13, p4o13_valid, p11i1_received, p11o0, p11o0_valid, p11o0_received, p11o1, p11o1_valid, p11o1_received);
	a12 a12_inst(clk, reset, p4o14, p4o14_valid, p12i0_received, p4o15, p4o15_valid, p12i1_received, p12o0, p12o0_valid, p12o0_received, p12o1, p12o1_valid, p12o1_received);
	a13 a13_inst(clk, reset, p4o8, p4o8_valid, p13i0_received, p4o9, p4o9_valid, p13i1_received, p13o0, p13o0_valid, p13o0_received, p13o1, p13o1_valid, p13o1_received);
	a14 a14_inst(clk, reset, p4o10, p4o10_valid, p14i0_received, p4o11, p4o11_valid, p14i1_received, p14o0, p14o0_valid, p14o0_received, p14o1, p14o1_valid, p14o1_received);
	a15 a15_inst(clk, reset, p4o12, p4o12_valid, p15i0_received, p4o13, p4o13_valid, p15i1_received, p15o0, p15o0_valid, p15o0_received, p15o1, p15o1_valid, p15o1_received);
	a16 a16_inst(clk, reset, p4o14, p4o14_valid, p16i0_received, p4o15, p4o15_valid, p16i1_received, p16o0, p16o0_valid, p16o0_received, p16o1, p16o1_valid, p16o1_received);
	a17 a17_inst(clk, reset, p4o8, p4o8_valid, p17i0_received, p4o9, p4o9_valid, p17i1_received, p17o0, p17o0_valid, p17o0_received, p17o1, p17o1_valid, p17o1_received);
	a18 a18_inst(clk, reset, p4o10, p4o10_valid, p18i0_received, p4o11, p4o11_valid, p18i1_received, p18o0, p18o0_valid, p18o0_received, p18o1, p18o1_valid, p18o1_received);
	a19 a19_inst(clk, reset, p4o12, p4o12_valid, p19i0_received, p4o13, p4o13_valid, p19i1_received, p19o0, p19o0_valid, p19o0_received, p19o1, p19o1_valid, p19o1_received);
	a20 a20_inst(clk, reset, p4o14, p4o14_valid, p20i0_received, p4o15, p4o15_valid, p20i1_received, p20o0, p20o0_valid, p20o0_received, p20o1, p20o1_valid, p20o1_received);

	assign o0 = p4o0;
	assign o0_valid = p4o0_valid;
	assign o1 = p4o1;
	assign o1_valid = p4o1_valid;
	assign o2 = p4o2;
	assign o2_valid = p4o2_valid;
	assign o3 = p4o3;
	assign o3_valid = p4o3_valid;
	assign o4 = p4o4;
	assign o4_valid = p4o4_valid;
	assign o5 = p4o5;
	assign o5_valid = p4o5_valid;
	assign o6 = p4o6;
	assign o6_valid = p4o6_valid;
	assign o7 = p4o7;
	assign o7_valid = p4o7_valid;

	assign p0o0_received = p4i8_received;
	assign p0o1_received = p4i9_received;
	assign p1o0_received = p4i10_received;
	assign p1o1_received = p4i11_received;
	assign p2o0_received = p4i12_received;
	assign p2o1_received = p4i13_received;
	assign p3o0_received = p4i14_received;
	assign p3o1_received = p4i15_received;
	assign p4o0_received = o0_received;
	assign p4o1_received = o1_received;
	assign p4o2_received = o2_received;
	assign p4o3_received = o3_received;
	assign p4o4_received = o4_received;
	assign p4o5_received = o5_received;
	assign p4o6_received = o6_received;
	assign p4o7_received = o7_received;
	assign p4o8_received = ( 1'b1 
		& (p5i0_received) 
		& (p9i0_received) 
		& (p13i0_received) 
		& (p17i0_received) 
		);
	assign p4o9_received = ( 1'b1 
		& (p5i1_received) 
		& (p9i1_received) 
		& (p13i1_received) 
		& (p17i1_received) 
		);
	assign p4o10_received = ( 1'b1 
		& (p6i0_received) 
		& (p10i0_received) 
		& (p14i0_received) 
		& (p18i0_received) 
		);
	assign p4o11_received = ( 1'b1 
		& (p6i1_received) 
		& (p10i1_received) 
		& (p14i1_received) 
		& (p18i1_received) 
		);
	assign p4o12_received = ( 1'b1 
		& (p7i0_received) 
		& (p11i0_received) 
		& (p15i0_received) 
		& (p19i0_received) 
		);
	assign p4o13_received = ( 1'b1 
		& (p7i1_received) 
		& (p11i1_received) 
		& (p15i1_received) 
		& (p19i1_received) 
		);
	assign p4o14_received = ( 1'b1 
		& (p8i0_received) 
		& (p12i0_received) 
		& (p16i0_received) 
		& (p20i0_received) 
		);
	assign p4o15_received = ( 1'b1 
		& (p8i1_received) 
		& (p12i1_received) 
		& (p16i1_received) 
		& (p20i1_received) 
		);
	assign p5o0_received = p0i0_received;
	assign p5o1_received = p0i1_received;
	assign p6o0_received = p0i2_received;
	assign p6o1_received = p0i3_received;
	assign p7o0_received = p0i4_received;
	assign p7o1_received = p0i5_received;
	assign p8o0_received = p0i6_received;
	assign p8o1_received = p0i7_received;
	assign p9o0_received = p1i0_received;
	assign p9o1_received = p1i1_received;
	assign p10o0_received = p1i2_received;
	assign p10o1_received = p1i3_received;
	assign p11o0_received = p1i4_received;
	assign p11o1_received = p1i5_received;
	assign p12o0_received = p1i6_received;
	assign p12o1_received = p1i7_received;
	assign p13o0_received = p2i0_received;
	assign p13o1_received = p2i1_received;
	assign p14o0_received = p2i2_received;
	assign p14o1_received = p2i3_received;
	assign p15o0_received = p2i4_received;
	assign p15o1_received = p2i5_received;
	assign p16o0_received = p2i6_received;
	assign p16o1_received = p2i7_received;
	assign p17o0_received = p3i0_received;
	assign p17o1_received = p3i1_received;
	assign p18o0_received = p3i2_received;
	assign p18o1_received = p3i3_received;
	assign p19o0_received = p3i4_received;
	assign p19o1_received = p3i5_received;
	assign p20o0_received = p3i6_received;
	assign p20o1_received = p3i7_received;
	assign i0_received = p4i0_received;
	assign i1_received = p4i1_received;
	assign i2_received = p4i2_received;
	assign i3_received = p4i3_received;
	assign i4_received = p4i4_received;
	assign i5_received = p4i5_received;
	assign i6_received = p4i6_received;
	assign i7_received = p4i7_received;

endmodule
`timescale 1ns/1ps
module p0rom(input [4:0] rom_bus, output [7:0] rom_value);
	reg [7:0] _rom [0:31];
	initial
	begin
	_rom[0] = 8'b00100000;
	_rom[1] = 8'b00101000;
	_rom[2] = 8'b01010000;
	_rom[3] = 8'b01011001;
	_rom[4] = 8'b00000100;
	_rom[5] = 8'b00001110;
	_rom[6] = 8'b01010010;
	_rom[7] = 8'b01011011;
	_rom[8] = 8'b00000100;
	_rom[9] = 8'b00001110;
	_rom[10] = 8'b01010100;
	_rom[11] = 8'b01011101;
	_rom[12] = 8'b00000100;
	_rom[13] = 8'b00001110;
	_rom[14] = 8'b01010110;
	_rom[15] = 8'b01011111;
	_rom[16] = 8'b00000100;
	_rom[17] = 8'b00001110;
	_rom[18] = 8'b10000000;
	_rom[19] = 8'b10001100;
	_rom[20] = 8'b01100000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p0(clock_signal, reset_signal, rom_bus, rom_value, i0, i0_valid, i0_received, i1, i1_valid, i1_received, i2, i2_valid, i2_received, i3, i3_valid, i3_received, i4, i4_valid, i4_received, i5, i5_valid, i5_received, i6, i6_valid, i6_received, i7, i7_valid, i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [7:0] rom_value;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=3'b000,          // Register addf
			CLR=3'b001,          // Clear register
			I2RW=3'b010,          // Input to register
			J=3'b011,          // Jump to a program location
			R2OWA=3'b100;          // Register to output

	localparam	R0=2'b00,		// Registers in the intructions
			R1=2'b01,
			R2=2'b10,
			R3=2'b11;
	localparam			I0=3'b000,
			I1=3'b001,
			I2=3'b010,
			I3=3'b011,
			I4=3'b100,
			I5=3'b101,
			I6=3'b110,
			I7=3'b111;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:0];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;

	wire [7:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_0_input_a;
	reg [31:0] adder_0_input_b;
	reg adder_0_input_a_stb;
	reg adder_0_input_b_stb;
	reg adder_0_output_z_ack;

	wire [31:0] adder_0_output_z;
	wire adder_0_output_z_stb;
	wire adder_0_input_a_ack;
	wire adder_0_input_b_ack;

	reg	[1:0] adder_0_state;
parameter adder_0_put_a         = 2'd0,
          adder_0_put_b         = 2'd1,
          adder_0_get_z         = 2'd2;
	adder_0 adder_0_inst (adder_0_input_a, adder_0_input_b, adder_0_input_a_stb, adder_0_input_b_stb, adder_0_output_z_ack, clock_signal, reset_signal, adder_0_output_z, adder_0_output_z_stb, adder_0_input_a_ack, adder_0_input_b_ack);


// Start of the component "header" for the opcode clr


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;
	reg i2_recv;
	reg i3_recv;
	reg i4_recv;
	reg i5_recv;
	reg i6_recv;
	reg i7_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i2_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I2 : begin
						if (i2_valid)
						begin
							i2_recv <= #1 1'b1;
						end else begin
							i2_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i2_valid)
						begin
							i2_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i2_valid)
					begin
						i2_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i3_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I3 : begin
						if (i3_valid)
						begin
							i3_recv <= #1 1'b1;
						end else begin
							i3_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i3_valid)
						begin
							i3_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i3_valid)
					begin
						i3_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i4_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I4 : begin
						if (i4_valid)
						begin
							i4_recv <= #1 1'b1;
						end else begin
							i4_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i4_valid)
						begin
							i4_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i4_valid)
					begin
						i4_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i5_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I5 : begin
						if (i5_valid)
						begin
							i5_recv <= #1 1'b1;
						end else begin
							i5_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i5_valid)
						begin
							i5_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i5_valid)
					begin
						i5_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i6_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I6 : begin
						if (i6_valid)
						begin
							i6_recv <= #1 1'b1;
						end else begin
							i6_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i6_valid)
						begin
							i6_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i6_valid)
					begin
						i6_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i7_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I7 : begin
						if (i7_valid)
						begin
							i7_recv <= #1 1'b1;
						end else begin
							i7_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i7_valid)
						begin
							i7_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i7_valid)
					begin
						i7_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				R2OWA: begin
					case (current_instruction[2])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				R2OWA: begin
					case (current_instruction[2])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode clr


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode r2owa

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b ", _r0, _r1, _r2, _r3);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode clr


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode r2owa


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode clr


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode r2owa

				case(current_instruction[7:5])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2:1])
							R2 : begin
							case (adder_0_state)
							adder_0_put_a : begin
								if (adder_0_input_a_ack) begin
									adder_0_input_a <= #1 _r0;
									adder_0_input_a_stb <= #1 1;
									adder_0_output_z_ack <= #1 0;
									adder_0_state <= #1 adder_0_put_b;
								end
							end
							adder_0_put_b : begin
								if (adder_0_input_b_ack) begin
									adder_0_input_b <= #1 _r2;
									adder_0_input_b_stb <= #1 1;
									adder_0_output_z_ack <= #1 0;
									adder_0_state <= #1 adder_0_get_z;
									adder_0_input_a_stb <= #1 0;
								end
							end
							adder_0_get_z : begin
								if (adder_0_output_z_stb) begin
									_r0 <= #1 adder_0_output_z;
									adder_0_output_z_ack <= #1 1;
									adder_0_state <= #1 adder_0_put_a;
									adder_0_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R2");
							end
							R3 : begin
							case (adder_0_state)
							adder_0_put_a : begin
								if (adder_0_input_a_ack) begin
									adder_0_input_a <= #1 _r0;
									adder_0_input_a_stb <= #1 1;
									adder_0_output_z_ack <= #1 0;
									adder_0_state <= #1 adder_0_put_b;
								end
							end
							adder_0_put_b : begin
								if (adder_0_input_b_ack) begin
									adder_0_input_b <= #1 _r3;
									adder_0_input_b_stb <= #1 1;
									adder_0_output_z_ack <= #1 0;
									adder_0_state <= #1 adder_0_get_z;
									adder_0_input_a_stb <= #1 0;
								end
							end
							adder_0_get_z : begin
								if (adder_0_output_z_stb) begin
									_r0 <= #1 adder_0_output_z;
									adder_0_output_z_ack <= #1 1;
									adder_0_state <= #1 adder_0_put_a;
									adder_0_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2:1])
							R2 : begin
							case (adder_0_state)
							adder_0_put_a : begin
								if (adder_0_input_a_ack) begin
									adder_0_input_a <= #1 _r1;
									adder_0_input_a_stb <= #1 1;
									adder_0_output_z_ack <= #1 0;
									adder_0_state <= #1 adder_0_put_b;
								end
							end
							adder_0_put_b : begin
								if (adder_0_input_b_ack) begin
									adder_0_input_b <= #1 _r2;
									adder_0_input_b_stb <= #1 1;
									adder_0_output_z_ack <= #1 0;
									adder_0_state <= #1 adder_0_get_z;
									adder_0_input_a_stb <= #1 0;
								end
							end
							adder_0_get_z : begin
								if (adder_0_output_z_stb) begin
									_r1 <= #1 adder_0_output_z;
									adder_0_output_z_ack <= #1 1;
									adder_0_state <= #1 adder_0_put_a;
									adder_0_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R1 R2");
							end
							R3 : begin
							case (adder_0_state)
							adder_0_put_a : begin
								if (adder_0_input_a_ack) begin
									adder_0_input_a <= #1 _r1;
									adder_0_input_a_stb <= #1 1;
									adder_0_output_z_ack <= #1 0;
									adder_0_state <= #1 adder_0_put_b;
								end
							end
							adder_0_put_b : begin
								if (adder_0_input_b_ack) begin
									adder_0_input_b <= #1 _r3;
									adder_0_input_b_stb <= #1 1;
									adder_0_output_z_ack <= #1 0;
									adder_0_state <= #1 adder_0_get_z;
									adder_0_input_a_stb <= #1 0;
								end
							end
							adder_0_get_z : begin
								if (adder_0_output_z_stb) begin
									_r1 <= #1 adder_0_output_z;
									adder_0_output_z_ack <= #1 1;
									adder_0_state <= #1 adder_0_put_a;
									adder_0_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R1 R3");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode clr

					CLR: begin
						case (current_instruction[4:3])
						R0 : begin
							_r0 <= #1 'b0;
							$display("CLR R0");
						end
						R1 : begin
							_r1 <= #1 'b0;
							$display("CLR R1");
						end
						R2 : begin
							_r2 <= #1 'b0;
							$display("CLR R2");
						end
						R3 : begin
							_r3 <= #1 'b0;
							$display("CLR R3");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r0 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r0 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r0 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r0 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r0 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r0 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I7");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r1 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r1 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r1 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r1 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r1 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r1 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I7");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r2 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r2 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r2 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r2 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r2 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r2 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I7");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r3 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r3 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r3 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r3 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r3 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r3 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I7");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[4:0];
						$display("J ", current_instruction[4:0]);
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						endcase
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign i2_received = i2_recv;
	assign i3_received = i3_recv;
	assign i4_received = i4_recv;
	assign i5_received = i5_recv;
	assign i6_received = i6_recv;
	assign i7_received = i7_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_0 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p10ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00111111001101010000010011110011;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00111111100000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p10rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p10(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_10_input_a;
	reg [31:0] adder_10_input_b;
	reg adder_10_input_a_stb;
	reg adder_10_input_b_stb;
	reg adder_10_output_z_ack;

	wire [31:0] adder_10_output_z;
	wire adder_10_output_z_stb;
	wire adder_10_input_a_ack;
	wire adder_10_input_b_ack;

	reg	[1:0] adder_10_state;
parameter adder_10_put_a         = 2'd0,
          adder_10_put_b         = 2'd1,
          adder_10_get_z         = 2'd2;
	adder_10 adder_10_inst (adder_10_input_a, adder_10_input_b, adder_10_input_a_stb, adder_10_input_b_stb, adder_10_output_z_ack, clock_signal, reset_signal, adder_10_output_z, adder_10_output_z_stb, adder_10_input_a_ack, adder_10_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_10_input_a;
	reg [31:0] multiplier_10_input_b;
	reg multiplier_10_input_a_stb;
	reg multiplier_10_input_b_stb;
	reg multiplier_10_output_z_ack;

	wire [31:0] multiplier_10_output_z;
	wire multiplier_10_output_z_stb;
	wire multiplier_10_input_a_ack;
	wire multiplier_10_input_b_ack;

	reg	[1:0] multiplier_10_state;
parameter multiplier_10_put_a         = 2'd0,
          multiplier_10_put_b         = 2'd1,
          multiplier_10_get_z         = 2'd2;
	multiplier_10 multiplier_10_inst (multiplier_10_input_a, multiplier_10_input_b, multiplier_10_input_a_stb, multiplier_10_input_b_stb, multiplier_10_output_z_ack, clock_signal, reset_signal, multiplier_10_output_z, multiplier_10_output_z_stb, multiplier_10_input_a_ack, multiplier_10_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_10_state)
							adder_10_put_a : begin
								if (adder_10_input_a_ack) begin
									adder_10_input_a <= #1 _r0;
									adder_10_input_a_stb <= #1 1;
									adder_10_output_z_ack <= #1 0;
									adder_10_state <= #1 adder_10_put_b;
								end
							end
							adder_10_put_b : begin
								if (adder_10_input_b_ack) begin
									adder_10_input_b <= #1 _r7;
									adder_10_input_b_stb <= #1 1;
									adder_10_output_z_ack <= #1 0;
									adder_10_state <= #1 adder_10_get_z;
									adder_10_input_a_stb <= #1 0;
								end
							end
							adder_10_get_z : begin
								if (adder_10_output_z_stb) begin
									_r0 <= #1 adder_10_output_z;
									adder_10_output_z_ack <= #1 1;
									adder_10_state <= #1 adder_10_put_a;
									adder_10_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_10_state)
							adder_10_put_a : begin
								if (adder_10_input_a_ack) begin
									adder_10_input_a <= #1 _r6;
									adder_10_input_a_stb <= #1 1;
									adder_10_output_z_ack <= #1 0;
									adder_10_state <= #1 adder_10_put_b;
								end
							end
							adder_10_put_b : begin
								if (adder_10_input_b_ack) begin
									adder_10_input_b <= #1 _r7;
									adder_10_input_b_stb <= #1 1;
									adder_10_output_z_ack <= #1 0;
									adder_10_state <= #1 adder_10_get_z;
									adder_10_input_a_stb <= #1 0;
								end
							end
							adder_10_get_z : begin
								if (adder_10_output_z_stb) begin
									_r6 <= #1 adder_10_output_z;
									adder_10_output_z_ack <= #1 1;
									adder_10_state <= #1 adder_10_put_a;
									adder_10_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_10_state)
							multiplier_10_put_a : begin
								if (multiplier_10_input_a_ack) begin
									multiplier_10_input_a <= #1 _r0;
									multiplier_10_input_a_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_put_b;
								end
							end
							multiplier_10_put_b : begin
								if (multiplier_10_input_b_ack) begin
									multiplier_10_input_b <= #1 _r3;
									multiplier_10_input_b_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_get_z;
									multiplier_10_input_a_stb <= #1 0;
								end
							end
							multiplier_10_get_z : begin
								if (multiplier_10_output_z_stb) begin
									_r0 <= #1 multiplier_10_output_z;
									multiplier_10_output_z_ack <= #1 1;
									multiplier_10_state <= #1 multiplier_10_put_a;
									multiplier_10_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_10_state)
							multiplier_10_put_a : begin
								if (multiplier_10_input_a_ack) begin
									multiplier_10_input_a <= #1 _r0;
									multiplier_10_input_a_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_put_b;
								end
							end
							multiplier_10_put_b : begin
								if (multiplier_10_input_b_ack) begin
									multiplier_10_input_b <= #1 _r4;
									multiplier_10_input_b_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_get_z;
									multiplier_10_input_a_stb <= #1 0;
								end
							end
							multiplier_10_get_z : begin
								if (multiplier_10_output_z_stb) begin
									_r0 <= #1 multiplier_10_output_z;
									multiplier_10_output_z_ack <= #1 1;
									multiplier_10_state <= #1 multiplier_10_put_a;
									multiplier_10_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_10_state)
							multiplier_10_put_a : begin
								if (multiplier_10_input_a_ack) begin
									multiplier_10_input_a <= #1 _r0;
									multiplier_10_input_a_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_put_b;
								end
							end
							multiplier_10_put_b : begin
								if (multiplier_10_input_b_ack) begin
									multiplier_10_input_b <= #1 _r5;
									multiplier_10_input_b_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_get_z;
									multiplier_10_input_a_stb <= #1 0;
								end
							end
							multiplier_10_get_z : begin
								if (multiplier_10_output_z_stb) begin
									_r0 <= #1 multiplier_10_output_z;
									multiplier_10_output_z_ack <= #1 1;
									multiplier_10_state <= #1 multiplier_10_put_a;
									multiplier_10_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_10_state)
							multiplier_10_put_a : begin
								if (multiplier_10_input_a_ack) begin
									multiplier_10_input_a <= #1 _r7;
									multiplier_10_input_a_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_put_b;
								end
							end
							multiplier_10_put_b : begin
								if (multiplier_10_input_b_ack) begin
									multiplier_10_input_b <= #1 _r3;
									multiplier_10_input_b_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_get_z;
									multiplier_10_input_a_stb <= #1 0;
								end
							end
							multiplier_10_get_z : begin
								if (multiplier_10_output_z_stb) begin
									_r7 <= #1 multiplier_10_output_z;
									multiplier_10_output_z_ack <= #1 1;
									multiplier_10_state <= #1 multiplier_10_put_a;
									multiplier_10_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_10_state)
							multiplier_10_put_a : begin
								if (multiplier_10_input_a_ack) begin
									multiplier_10_input_a <= #1 _r7;
									multiplier_10_input_a_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_put_b;
								end
							end
							multiplier_10_put_b : begin
								if (multiplier_10_input_b_ack) begin
									multiplier_10_input_b <= #1 _r4;
									multiplier_10_input_b_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_get_z;
									multiplier_10_input_a_stb <= #1 0;
								end
							end
							multiplier_10_get_z : begin
								if (multiplier_10_output_z_stb) begin
									_r7 <= #1 multiplier_10_output_z;
									multiplier_10_output_z_ack <= #1 1;
									multiplier_10_state <= #1 multiplier_10_put_a;
									multiplier_10_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_10_state)
							multiplier_10_put_a : begin
								if (multiplier_10_input_a_ack) begin
									multiplier_10_input_a <= #1 _r7;
									multiplier_10_input_a_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_put_b;
								end
							end
							multiplier_10_put_b : begin
								if (multiplier_10_input_b_ack) begin
									multiplier_10_input_b <= #1 _r5;
									multiplier_10_input_b_stb <= #1 1;
									multiplier_10_output_z_ack <= #1 0;
									multiplier_10_state <= #1 multiplier_10_get_z;
									multiplier_10_input_a_stb <= #1 0;
								end
							end
							multiplier_10_get_z : begin
								if (multiplier_10_output_z_stb) begin
									_r7 <= #1 multiplier_10_output_z;
									multiplier_10_output_z_ack <= #1 1;
									multiplier_10_state <= #1 multiplier_10_put_a;
									multiplier_10_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_10 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_10 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p11ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00000000000000000000000000000000;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p11rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p11(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_11_input_a;
	reg [31:0] adder_11_input_b;
	reg adder_11_input_a_stb;
	reg adder_11_input_b_stb;
	reg adder_11_output_z_ack;

	wire [31:0] adder_11_output_z;
	wire adder_11_output_z_stb;
	wire adder_11_input_a_ack;
	wire adder_11_input_b_ack;

	reg	[1:0] adder_11_state;
parameter adder_11_put_a         = 2'd0,
          adder_11_put_b         = 2'd1,
          adder_11_get_z         = 2'd2;
	adder_11 adder_11_inst (adder_11_input_a, adder_11_input_b, adder_11_input_a_stb, adder_11_input_b_stb, adder_11_output_z_ack, clock_signal, reset_signal, adder_11_output_z, adder_11_output_z_stb, adder_11_input_a_ack, adder_11_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_11_input_a;
	reg [31:0] multiplier_11_input_b;
	reg multiplier_11_input_a_stb;
	reg multiplier_11_input_b_stb;
	reg multiplier_11_output_z_ack;

	wire [31:0] multiplier_11_output_z;
	wire multiplier_11_output_z_stb;
	wire multiplier_11_input_a_ack;
	wire multiplier_11_input_b_ack;

	reg	[1:0] multiplier_11_state;
parameter multiplier_11_put_a         = 2'd0,
          multiplier_11_put_b         = 2'd1,
          multiplier_11_get_z         = 2'd2;
	multiplier_11 multiplier_11_inst (multiplier_11_input_a, multiplier_11_input_b, multiplier_11_input_a_stb, multiplier_11_input_b_stb, multiplier_11_output_z_ack, clock_signal, reset_signal, multiplier_11_output_z, multiplier_11_output_z_stb, multiplier_11_input_a_ack, multiplier_11_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_11_state)
							adder_11_put_a : begin
								if (adder_11_input_a_ack) begin
									adder_11_input_a <= #1 _r0;
									adder_11_input_a_stb <= #1 1;
									adder_11_output_z_ack <= #1 0;
									adder_11_state <= #1 adder_11_put_b;
								end
							end
							adder_11_put_b : begin
								if (adder_11_input_b_ack) begin
									adder_11_input_b <= #1 _r7;
									adder_11_input_b_stb <= #1 1;
									adder_11_output_z_ack <= #1 0;
									adder_11_state <= #1 adder_11_get_z;
									adder_11_input_a_stb <= #1 0;
								end
							end
							adder_11_get_z : begin
								if (adder_11_output_z_stb) begin
									_r0 <= #1 adder_11_output_z;
									adder_11_output_z_ack <= #1 1;
									adder_11_state <= #1 adder_11_put_a;
									adder_11_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_11_state)
							adder_11_put_a : begin
								if (adder_11_input_a_ack) begin
									adder_11_input_a <= #1 _r6;
									adder_11_input_a_stb <= #1 1;
									adder_11_output_z_ack <= #1 0;
									adder_11_state <= #1 adder_11_put_b;
								end
							end
							adder_11_put_b : begin
								if (adder_11_input_b_ack) begin
									adder_11_input_b <= #1 _r7;
									adder_11_input_b_stb <= #1 1;
									adder_11_output_z_ack <= #1 0;
									adder_11_state <= #1 adder_11_get_z;
									adder_11_input_a_stb <= #1 0;
								end
							end
							adder_11_get_z : begin
								if (adder_11_output_z_stb) begin
									_r6 <= #1 adder_11_output_z;
									adder_11_output_z_ack <= #1 1;
									adder_11_state <= #1 adder_11_put_a;
									adder_11_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_11_state)
							multiplier_11_put_a : begin
								if (multiplier_11_input_a_ack) begin
									multiplier_11_input_a <= #1 _r0;
									multiplier_11_input_a_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_put_b;
								end
							end
							multiplier_11_put_b : begin
								if (multiplier_11_input_b_ack) begin
									multiplier_11_input_b <= #1 _r3;
									multiplier_11_input_b_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_get_z;
									multiplier_11_input_a_stb <= #1 0;
								end
							end
							multiplier_11_get_z : begin
								if (multiplier_11_output_z_stb) begin
									_r0 <= #1 multiplier_11_output_z;
									multiplier_11_output_z_ack <= #1 1;
									multiplier_11_state <= #1 multiplier_11_put_a;
									multiplier_11_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_11_state)
							multiplier_11_put_a : begin
								if (multiplier_11_input_a_ack) begin
									multiplier_11_input_a <= #1 _r0;
									multiplier_11_input_a_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_put_b;
								end
							end
							multiplier_11_put_b : begin
								if (multiplier_11_input_b_ack) begin
									multiplier_11_input_b <= #1 _r4;
									multiplier_11_input_b_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_get_z;
									multiplier_11_input_a_stb <= #1 0;
								end
							end
							multiplier_11_get_z : begin
								if (multiplier_11_output_z_stb) begin
									_r0 <= #1 multiplier_11_output_z;
									multiplier_11_output_z_ack <= #1 1;
									multiplier_11_state <= #1 multiplier_11_put_a;
									multiplier_11_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_11_state)
							multiplier_11_put_a : begin
								if (multiplier_11_input_a_ack) begin
									multiplier_11_input_a <= #1 _r0;
									multiplier_11_input_a_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_put_b;
								end
							end
							multiplier_11_put_b : begin
								if (multiplier_11_input_b_ack) begin
									multiplier_11_input_b <= #1 _r5;
									multiplier_11_input_b_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_get_z;
									multiplier_11_input_a_stb <= #1 0;
								end
							end
							multiplier_11_get_z : begin
								if (multiplier_11_output_z_stb) begin
									_r0 <= #1 multiplier_11_output_z;
									multiplier_11_output_z_ack <= #1 1;
									multiplier_11_state <= #1 multiplier_11_put_a;
									multiplier_11_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_11_state)
							multiplier_11_put_a : begin
								if (multiplier_11_input_a_ack) begin
									multiplier_11_input_a <= #1 _r7;
									multiplier_11_input_a_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_put_b;
								end
							end
							multiplier_11_put_b : begin
								if (multiplier_11_input_b_ack) begin
									multiplier_11_input_b <= #1 _r3;
									multiplier_11_input_b_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_get_z;
									multiplier_11_input_a_stb <= #1 0;
								end
							end
							multiplier_11_get_z : begin
								if (multiplier_11_output_z_stb) begin
									_r7 <= #1 multiplier_11_output_z;
									multiplier_11_output_z_ack <= #1 1;
									multiplier_11_state <= #1 multiplier_11_put_a;
									multiplier_11_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_11_state)
							multiplier_11_put_a : begin
								if (multiplier_11_input_a_ack) begin
									multiplier_11_input_a <= #1 _r7;
									multiplier_11_input_a_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_put_b;
								end
							end
							multiplier_11_put_b : begin
								if (multiplier_11_input_b_ack) begin
									multiplier_11_input_b <= #1 _r4;
									multiplier_11_input_b_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_get_z;
									multiplier_11_input_a_stb <= #1 0;
								end
							end
							multiplier_11_get_z : begin
								if (multiplier_11_output_z_stb) begin
									_r7 <= #1 multiplier_11_output_z;
									multiplier_11_output_z_ack <= #1 1;
									multiplier_11_state <= #1 multiplier_11_put_a;
									multiplier_11_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_11_state)
							multiplier_11_put_a : begin
								if (multiplier_11_input_a_ack) begin
									multiplier_11_input_a <= #1 _r7;
									multiplier_11_input_a_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_put_b;
								end
							end
							multiplier_11_put_b : begin
								if (multiplier_11_input_b_ack) begin
									multiplier_11_input_b <= #1 _r5;
									multiplier_11_input_b_stb <= #1 1;
									multiplier_11_output_z_ack <= #1 0;
									multiplier_11_state <= #1 multiplier_11_get_z;
									multiplier_11_input_a_stb <= #1 0;
								end
							end
							multiplier_11_get_z : begin
								if (multiplier_11_output_z_stb) begin
									_r7 <= #1 multiplier_11_output_z;
									multiplier_11_output_z_ack <= #1 1;
									multiplier_11_state <= #1 multiplier_11_put_a;
									multiplier_11_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_11 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_11 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p12ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00111111001101010000010011110011;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p12rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p12(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_12_input_a;
	reg [31:0] adder_12_input_b;
	reg adder_12_input_a_stb;
	reg adder_12_input_b_stb;
	reg adder_12_output_z_ack;

	wire [31:0] adder_12_output_z;
	wire adder_12_output_z_stb;
	wire adder_12_input_a_ack;
	wire adder_12_input_b_ack;

	reg	[1:0] adder_12_state;
parameter adder_12_put_a         = 2'd0,
          adder_12_put_b         = 2'd1,
          adder_12_get_z         = 2'd2;
	adder_12 adder_12_inst (adder_12_input_a, adder_12_input_b, adder_12_input_a_stb, adder_12_input_b_stb, adder_12_output_z_ack, clock_signal, reset_signal, adder_12_output_z, adder_12_output_z_stb, adder_12_input_a_ack, adder_12_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_12_input_a;
	reg [31:0] multiplier_12_input_b;
	reg multiplier_12_input_a_stb;
	reg multiplier_12_input_b_stb;
	reg multiplier_12_output_z_ack;

	wire [31:0] multiplier_12_output_z;
	wire multiplier_12_output_z_stb;
	wire multiplier_12_input_a_ack;
	wire multiplier_12_input_b_ack;

	reg	[1:0] multiplier_12_state;
parameter multiplier_12_put_a         = 2'd0,
          multiplier_12_put_b         = 2'd1,
          multiplier_12_get_z         = 2'd2;
	multiplier_12 multiplier_12_inst (multiplier_12_input_a, multiplier_12_input_b, multiplier_12_input_a_stb, multiplier_12_input_b_stb, multiplier_12_output_z_ack, clock_signal, reset_signal, multiplier_12_output_z, multiplier_12_output_z_stb, multiplier_12_input_a_ack, multiplier_12_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_12_state)
							adder_12_put_a : begin
								if (adder_12_input_a_ack) begin
									adder_12_input_a <= #1 _r0;
									adder_12_input_a_stb <= #1 1;
									adder_12_output_z_ack <= #1 0;
									adder_12_state <= #1 adder_12_put_b;
								end
							end
							adder_12_put_b : begin
								if (adder_12_input_b_ack) begin
									adder_12_input_b <= #1 _r7;
									adder_12_input_b_stb <= #1 1;
									adder_12_output_z_ack <= #1 0;
									adder_12_state <= #1 adder_12_get_z;
									adder_12_input_a_stb <= #1 0;
								end
							end
							adder_12_get_z : begin
								if (adder_12_output_z_stb) begin
									_r0 <= #1 adder_12_output_z;
									adder_12_output_z_ack <= #1 1;
									adder_12_state <= #1 adder_12_put_a;
									adder_12_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_12_state)
							adder_12_put_a : begin
								if (adder_12_input_a_ack) begin
									adder_12_input_a <= #1 _r6;
									adder_12_input_a_stb <= #1 1;
									adder_12_output_z_ack <= #1 0;
									adder_12_state <= #1 adder_12_put_b;
								end
							end
							adder_12_put_b : begin
								if (adder_12_input_b_ack) begin
									adder_12_input_b <= #1 _r7;
									adder_12_input_b_stb <= #1 1;
									adder_12_output_z_ack <= #1 0;
									adder_12_state <= #1 adder_12_get_z;
									adder_12_input_a_stb <= #1 0;
								end
							end
							adder_12_get_z : begin
								if (adder_12_output_z_stb) begin
									_r6 <= #1 adder_12_output_z;
									adder_12_output_z_ack <= #1 1;
									adder_12_state <= #1 adder_12_put_a;
									adder_12_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_12_state)
							multiplier_12_put_a : begin
								if (multiplier_12_input_a_ack) begin
									multiplier_12_input_a <= #1 _r0;
									multiplier_12_input_a_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_put_b;
								end
							end
							multiplier_12_put_b : begin
								if (multiplier_12_input_b_ack) begin
									multiplier_12_input_b <= #1 _r3;
									multiplier_12_input_b_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_get_z;
									multiplier_12_input_a_stb <= #1 0;
								end
							end
							multiplier_12_get_z : begin
								if (multiplier_12_output_z_stb) begin
									_r0 <= #1 multiplier_12_output_z;
									multiplier_12_output_z_ack <= #1 1;
									multiplier_12_state <= #1 multiplier_12_put_a;
									multiplier_12_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_12_state)
							multiplier_12_put_a : begin
								if (multiplier_12_input_a_ack) begin
									multiplier_12_input_a <= #1 _r0;
									multiplier_12_input_a_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_put_b;
								end
							end
							multiplier_12_put_b : begin
								if (multiplier_12_input_b_ack) begin
									multiplier_12_input_b <= #1 _r4;
									multiplier_12_input_b_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_get_z;
									multiplier_12_input_a_stb <= #1 0;
								end
							end
							multiplier_12_get_z : begin
								if (multiplier_12_output_z_stb) begin
									_r0 <= #1 multiplier_12_output_z;
									multiplier_12_output_z_ack <= #1 1;
									multiplier_12_state <= #1 multiplier_12_put_a;
									multiplier_12_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_12_state)
							multiplier_12_put_a : begin
								if (multiplier_12_input_a_ack) begin
									multiplier_12_input_a <= #1 _r0;
									multiplier_12_input_a_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_put_b;
								end
							end
							multiplier_12_put_b : begin
								if (multiplier_12_input_b_ack) begin
									multiplier_12_input_b <= #1 _r5;
									multiplier_12_input_b_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_get_z;
									multiplier_12_input_a_stb <= #1 0;
								end
							end
							multiplier_12_get_z : begin
								if (multiplier_12_output_z_stb) begin
									_r0 <= #1 multiplier_12_output_z;
									multiplier_12_output_z_ack <= #1 1;
									multiplier_12_state <= #1 multiplier_12_put_a;
									multiplier_12_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_12_state)
							multiplier_12_put_a : begin
								if (multiplier_12_input_a_ack) begin
									multiplier_12_input_a <= #1 _r7;
									multiplier_12_input_a_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_put_b;
								end
							end
							multiplier_12_put_b : begin
								if (multiplier_12_input_b_ack) begin
									multiplier_12_input_b <= #1 _r3;
									multiplier_12_input_b_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_get_z;
									multiplier_12_input_a_stb <= #1 0;
								end
							end
							multiplier_12_get_z : begin
								if (multiplier_12_output_z_stb) begin
									_r7 <= #1 multiplier_12_output_z;
									multiplier_12_output_z_ack <= #1 1;
									multiplier_12_state <= #1 multiplier_12_put_a;
									multiplier_12_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_12_state)
							multiplier_12_put_a : begin
								if (multiplier_12_input_a_ack) begin
									multiplier_12_input_a <= #1 _r7;
									multiplier_12_input_a_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_put_b;
								end
							end
							multiplier_12_put_b : begin
								if (multiplier_12_input_b_ack) begin
									multiplier_12_input_b <= #1 _r4;
									multiplier_12_input_b_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_get_z;
									multiplier_12_input_a_stb <= #1 0;
								end
							end
							multiplier_12_get_z : begin
								if (multiplier_12_output_z_stb) begin
									_r7 <= #1 multiplier_12_output_z;
									multiplier_12_output_z_ack <= #1 1;
									multiplier_12_state <= #1 multiplier_12_put_a;
									multiplier_12_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_12_state)
							multiplier_12_put_a : begin
								if (multiplier_12_input_a_ack) begin
									multiplier_12_input_a <= #1 _r7;
									multiplier_12_input_a_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_put_b;
								end
							end
							multiplier_12_put_b : begin
								if (multiplier_12_input_b_ack) begin
									multiplier_12_input_b <= #1 _r5;
									multiplier_12_input_b_stb <= #1 1;
									multiplier_12_output_z_ack <= #1 0;
									multiplier_12_state <= #1 multiplier_12_get_z;
									multiplier_12_input_a_stb <= #1 0;
								end
							end
							multiplier_12_get_z : begin
								if (multiplier_12_output_z_stb) begin
									_r7 <= #1 multiplier_12_output_z;
									multiplier_12_output_z_ack <= #1 1;
									multiplier_12_state <= #1 multiplier_12_put_a;
									multiplier_12_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_12 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_12 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p13ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00111111001101010000010011110011;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p13rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p13(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_13_input_a;
	reg [31:0] adder_13_input_b;
	reg adder_13_input_a_stb;
	reg adder_13_input_b_stb;
	reg adder_13_output_z_ack;

	wire [31:0] adder_13_output_z;
	wire adder_13_output_z_stb;
	wire adder_13_input_a_ack;
	wire adder_13_input_b_ack;

	reg	[1:0] adder_13_state;
parameter adder_13_put_a         = 2'd0,
          adder_13_put_b         = 2'd1,
          adder_13_get_z         = 2'd2;
	adder_13 adder_13_inst (adder_13_input_a, adder_13_input_b, adder_13_input_a_stb, adder_13_input_b_stb, adder_13_output_z_ack, clock_signal, reset_signal, adder_13_output_z, adder_13_output_z_stb, adder_13_input_a_ack, adder_13_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_13_input_a;
	reg [31:0] multiplier_13_input_b;
	reg multiplier_13_input_a_stb;
	reg multiplier_13_input_b_stb;
	reg multiplier_13_output_z_ack;

	wire [31:0] multiplier_13_output_z;
	wire multiplier_13_output_z_stb;
	wire multiplier_13_input_a_ack;
	wire multiplier_13_input_b_ack;

	reg	[1:0] multiplier_13_state;
parameter multiplier_13_put_a         = 2'd0,
          multiplier_13_put_b         = 2'd1,
          multiplier_13_get_z         = 2'd2;
	multiplier_13 multiplier_13_inst (multiplier_13_input_a, multiplier_13_input_b, multiplier_13_input_a_stb, multiplier_13_input_b_stb, multiplier_13_output_z_ack, clock_signal, reset_signal, multiplier_13_output_z, multiplier_13_output_z_stb, multiplier_13_input_a_ack, multiplier_13_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_13_state)
							adder_13_put_a : begin
								if (adder_13_input_a_ack) begin
									adder_13_input_a <= #1 _r0;
									adder_13_input_a_stb <= #1 1;
									adder_13_output_z_ack <= #1 0;
									adder_13_state <= #1 adder_13_put_b;
								end
							end
							adder_13_put_b : begin
								if (adder_13_input_b_ack) begin
									adder_13_input_b <= #1 _r7;
									adder_13_input_b_stb <= #1 1;
									adder_13_output_z_ack <= #1 0;
									adder_13_state <= #1 adder_13_get_z;
									adder_13_input_a_stb <= #1 0;
								end
							end
							adder_13_get_z : begin
								if (adder_13_output_z_stb) begin
									_r0 <= #1 adder_13_output_z;
									adder_13_output_z_ack <= #1 1;
									adder_13_state <= #1 adder_13_put_a;
									adder_13_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_13_state)
							adder_13_put_a : begin
								if (adder_13_input_a_ack) begin
									adder_13_input_a <= #1 _r6;
									adder_13_input_a_stb <= #1 1;
									adder_13_output_z_ack <= #1 0;
									adder_13_state <= #1 adder_13_put_b;
								end
							end
							adder_13_put_b : begin
								if (adder_13_input_b_ack) begin
									adder_13_input_b <= #1 _r7;
									adder_13_input_b_stb <= #1 1;
									adder_13_output_z_ack <= #1 0;
									adder_13_state <= #1 adder_13_get_z;
									adder_13_input_a_stb <= #1 0;
								end
							end
							adder_13_get_z : begin
								if (adder_13_output_z_stb) begin
									_r6 <= #1 adder_13_output_z;
									adder_13_output_z_ack <= #1 1;
									adder_13_state <= #1 adder_13_put_a;
									adder_13_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_13_state)
							multiplier_13_put_a : begin
								if (multiplier_13_input_a_ack) begin
									multiplier_13_input_a <= #1 _r0;
									multiplier_13_input_a_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_put_b;
								end
							end
							multiplier_13_put_b : begin
								if (multiplier_13_input_b_ack) begin
									multiplier_13_input_b <= #1 _r3;
									multiplier_13_input_b_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_get_z;
									multiplier_13_input_a_stb <= #1 0;
								end
							end
							multiplier_13_get_z : begin
								if (multiplier_13_output_z_stb) begin
									_r0 <= #1 multiplier_13_output_z;
									multiplier_13_output_z_ack <= #1 1;
									multiplier_13_state <= #1 multiplier_13_put_a;
									multiplier_13_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_13_state)
							multiplier_13_put_a : begin
								if (multiplier_13_input_a_ack) begin
									multiplier_13_input_a <= #1 _r0;
									multiplier_13_input_a_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_put_b;
								end
							end
							multiplier_13_put_b : begin
								if (multiplier_13_input_b_ack) begin
									multiplier_13_input_b <= #1 _r4;
									multiplier_13_input_b_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_get_z;
									multiplier_13_input_a_stb <= #1 0;
								end
							end
							multiplier_13_get_z : begin
								if (multiplier_13_output_z_stb) begin
									_r0 <= #1 multiplier_13_output_z;
									multiplier_13_output_z_ack <= #1 1;
									multiplier_13_state <= #1 multiplier_13_put_a;
									multiplier_13_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_13_state)
							multiplier_13_put_a : begin
								if (multiplier_13_input_a_ack) begin
									multiplier_13_input_a <= #1 _r0;
									multiplier_13_input_a_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_put_b;
								end
							end
							multiplier_13_put_b : begin
								if (multiplier_13_input_b_ack) begin
									multiplier_13_input_b <= #1 _r5;
									multiplier_13_input_b_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_get_z;
									multiplier_13_input_a_stb <= #1 0;
								end
							end
							multiplier_13_get_z : begin
								if (multiplier_13_output_z_stb) begin
									_r0 <= #1 multiplier_13_output_z;
									multiplier_13_output_z_ack <= #1 1;
									multiplier_13_state <= #1 multiplier_13_put_a;
									multiplier_13_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_13_state)
							multiplier_13_put_a : begin
								if (multiplier_13_input_a_ack) begin
									multiplier_13_input_a <= #1 _r7;
									multiplier_13_input_a_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_put_b;
								end
							end
							multiplier_13_put_b : begin
								if (multiplier_13_input_b_ack) begin
									multiplier_13_input_b <= #1 _r3;
									multiplier_13_input_b_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_get_z;
									multiplier_13_input_a_stb <= #1 0;
								end
							end
							multiplier_13_get_z : begin
								if (multiplier_13_output_z_stb) begin
									_r7 <= #1 multiplier_13_output_z;
									multiplier_13_output_z_ack <= #1 1;
									multiplier_13_state <= #1 multiplier_13_put_a;
									multiplier_13_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_13_state)
							multiplier_13_put_a : begin
								if (multiplier_13_input_a_ack) begin
									multiplier_13_input_a <= #1 _r7;
									multiplier_13_input_a_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_put_b;
								end
							end
							multiplier_13_put_b : begin
								if (multiplier_13_input_b_ack) begin
									multiplier_13_input_b <= #1 _r4;
									multiplier_13_input_b_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_get_z;
									multiplier_13_input_a_stb <= #1 0;
								end
							end
							multiplier_13_get_z : begin
								if (multiplier_13_output_z_stb) begin
									_r7 <= #1 multiplier_13_output_z;
									multiplier_13_output_z_ack <= #1 1;
									multiplier_13_state <= #1 multiplier_13_put_a;
									multiplier_13_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_13_state)
							multiplier_13_put_a : begin
								if (multiplier_13_input_a_ack) begin
									multiplier_13_input_a <= #1 _r7;
									multiplier_13_input_a_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_put_b;
								end
							end
							multiplier_13_put_b : begin
								if (multiplier_13_input_b_ack) begin
									multiplier_13_input_b <= #1 _r5;
									multiplier_13_input_b_stb <= #1 1;
									multiplier_13_output_z_ack <= #1 0;
									multiplier_13_state <= #1 multiplier_13_get_z;
									multiplier_13_input_a_stb <= #1 0;
								end
							end
							multiplier_13_get_z : begin
								if (multiplier_13_output_z_stb) begin
									_r7 <= #1 multiplier_13_output_z;
									multiplier_13_output_z_ack <= #1 1;
									multiplier_13_state <= #1 multiplier_13_put_a;
									multiplier_13_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_13 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_13 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p14ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00000000000000000000000000000000;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p14rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p14(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_14_input_a;
	reg [31:0] adder_14_input_b;
	reg adder_14_input_a_stb;
	reg adder_14_input_b_stb;
	reg adder_14_output_z_ack;

	wire [31:0] adder_14_output_z;
	wire adder_14_output_z_stb;
	wire adder_14_input_a_ack;
	wire adder_14_input_b_ack;

	reg	[1:0] adder_14_state;
parameter adder_14_put_a         = 2'd0,
          adder_14_put_b         = 2'd1,
          adder_14_get_z         = 2'd2;
	adder_14 adder_14_inst (adder_14_input_a, adder_14_input_b, adder_14_input_a_stb, adder_14_input_b_stb, adder_14_output_z_ack, clock_signal, reset_signal, adder_14_output_z, adder_14_output_z_stb, adder_14_input_a_ack, adder_14_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_14_input_a;
	reg [31:0] multiplier_14_input_b;
	reg multiplier_14_input_a_stb;
	reg multiplier_14_input_b_stb;
	reg multiplier_14_output_z_ack;

	wire [31:0] multiplier_14_output_z;
	wire multiplier_14_output_z_stb;
	wire multiplier_14_input_a_ack;
	wire multiplier_14_input_b_ack;

	reg	[1:0] multiplier_14_state;
parameter multiplier_14_put_a         = 2'd0,
          multiplier_14_put_b         = 2'd1,
          multiplier_14_get_z         = 2'd2;
	multiplier_14 multiplier_14_inst (multiplier_14_input_a, multiplier_14_input_b, multiplier_14_input_a_stb, multiplier_14_input_b_stb, multiplier_14_output_z_ack, clock_signal, reset_signal, multiplier_14_output_z, multiplier_14_output_z_stb, multiplier_14_input_a_ack, multiplier_14_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_14_state)
							adder_14_put_a : begin
								if (adder_14_input_a_ack) begin
									adder_14_input_a <= #1 _r0;
									adder_14_input_a_stb <= #1 1;
									adder_14_output_z_ack <= #1 0;
									adder_14_state <= #1 adder_14_put_b;
								end
							end
							adder_14_put_b : begin
								if (adder_14_input_b_ack) begin
									adder_14_input_b <= #1 _r7;
									adder_14_input_b_stb <= #1 1;
									adder_14_output_z_ack <= #1 0;
									adder_14_state <= #1 adder_14_get_z;
									adder_14_input_a_stb <= #1 0;
								end
							end
							adder_14_get_z : begin
								if (adder_14_output_z_stb) begin
									_r0 <= #1 adder_14_output_z;
									adder_14_output_z_ack <= #1 1;
									adder_14_state <= #1 adder_14_put_a;
									adder_14_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_14_state)
							adder_14_put_a : begin
								if (adder_14_input_a_ack) begin
									adder_14_input_a <= #1 _r6;
									adder_14_input_a_stb <= #1 1;
									adder_14_output_z_ack <= #1 0;
									adder_14_state <= #1 adder_14_put_b;
								end
							end
							adder_14_put_b : begin
								if (adder_14_input_b_ack) begin
									adder_14_input_b <= #1 _r7;
									adder_14_input_b_stb <= #1 1;
									adder_14_output_z_ack <= #1 0;
									adder_14_state <= #1 adder_14_get_z;
									adder_14_input_a_stb <= #1 0;
								end
							end
							adder_14_get_z : begin
								if (adder_14_output_z_stb) begin
									_r6 <= #1 adder_14_output_z;
									adder_14_output_z_ack <= #1 1;
									adder_14_state <= #1 adder_14_put_a;
									adder_14_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_14_state)
							multiplier_14_put_a : begin
								if (multiplier_14_input_a_ack) begin
									multiplier_14_input_a <= #1 _r0;
									multiplier_14_input_a_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_put_b;
								end
							end
							multiplier_14_put_b : begin
								if (multiplier_14_input_b_ack) begin
									multiplier_14_input_b <= #1 _r3;
									multiplier_14_input_b_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_get_z;
									multiplier_14_input_a_stb <= #1 0;
								end
							end
							multiplier_14_get_z : begin
								if (multiplier_14_output_z_stb) begin
									_r0 <= #1 multiplier_14_output_z;
									multiplier_14_output_z_ack <= #1 1;
									multiplier_14_state <= #1 multiplier_14_put_a;
									multiplier_14_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_14_state)
							multiplier_14_put_a : begin
								if (multiplier_14_input_a_ack) begin
									multiplier_14_input_a <= #1 _r0;
									multiplier_14_input_a_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_put_b;
								end
							end
							multiplier_14_put_b : begin
								if (multiplier_14_input_b_ack) begin
									multiplier_14_input_b <= #1 _r4;
									multiplier_14_input_b_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_get_z;
									multiplier_14_input_a_stb <= #1 0;
								end
							end
							multiplier_14_get_z : begin
								if (multiplier_14_output_z_stb) begin
									_r0 <= #1 multiplier_14_output_z;
									multiplier_14_output_z_ack <= #1 1;
									multiplier_14_state <= #1 multiplier_14_put_a;
									multiplier_14_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_14_state)
							multiplier_14_put_a : begin
								if (multiplier_14_input_a_ack) begin
									multiplier_14_input_a <= #1 _r0;
									multiplier_14_input_a_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_put_b;
								end
							end
							multiplier_14_put_b : begin
								if (multiplier_14_input_b_ack) begin
									multiplier_14_input_b <= #1 _r5;
									multiplier_14_input_b_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_get_z;
									multiplier_14_input_a_stb <= #1 0;
								end
							end
							multiplier_14_get_z : begin
								if (multiplier_14_output_z_stb) begin
									_r0 <= #1 multiplier_14_output_z;
									multiplier_14_output_z_ack <= #1 1;
									multiplier_14_state <= #1 multiplier_14_put_a;
									multiplier_14_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_14_state)
							multiplier_14_put_a : begin
								if (multiplier_14_input_a_ack) begin
									multiplier_14_input_a <= #1 _r7;
									multiplier_14_input_a_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_put_b;
								end
							end
							multiplier_14_put_b : begin
								if (multiplier_14_input_b_ack) begin
									multiplier_14_input_b <= #1 _r3;
									multiplier_14_input_b_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_get_z;
									multiplier_14_input_a_stb <= #1 0;
								end
							end
							multiplier_14_get_z : begin
								if (multiplier_14_output_z_stb) begin
									_r7 <= #1 multiplier_14_output_z;
									multiplier_14_output_z_ack <= #1 1;
									multiplier_14_state <= #1 multiplier_14_put_a;
									multiplier_14_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_14_state)
							multiplier_14_put_a : begin
								if (multiplier_14_input_a_ack) begin
									multiplier_14_input_a <= #1 _r7;
									multiplier_14_input_a_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_put_b;
								end
							end
							multiplier_14_put_b : begin
								if (multiplier_14_input_b_ack) begin
									multiplier_14_input_b <= #1 _r4;
									multiplier_14_input_b_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_get_z;
									multiplier_14_input_a_stb <= #1 0;
								end
							end
							multiplier_14_get_z : begin
								if (multiplier_14_output_z_stb) begin
									_r7 <= #1 multiplier_14_output_z;
									multiplier_14_output_z_ack <= #1 1;
									multiplier_14_state <= #1 multiplier_14_put_a;
									multiplier_14_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_14_state)
							multiplier_14_put_a : begin
								if (multiplier_14_input_a_ack) begin
									multiplier_14_input_a <= #1 _r7;
									multiplier_14_input_a_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_put_b;
								end
							end
							multiplier_14_put_b : begin
								if (multiplier_14_input_b_ack) begin
									multiplier_14_input_b <= #1 _r5;
									multiplier_14_input_b_stb <= #1 1;
									multiplier_14_output_z_ack <= #1 0;
									multiplier_14_state <= #1 multiplier_14_get_z;
									multiplier_14_input_a_stb <= #1 0;
								end
							end
							multiplier_14_get_z : begin
								if (multiplier_14_output_z_stb) begin
									_r7 <= #1 multiplier_14_output_z;
									multiplier_14_output_z_ack <= #1 1;
									multiplier_14_state <= #1 multiplier_14_put_a;
									multiplier_14_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_14 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_14 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p15ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b10111111001101010000010011110011;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p15rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p15(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_15_input_a;
	reg [31:0] adder_15_input_b;
	reg adder_15_input_a_stb;
	reg adder_15_input_b_stb;
	reg adder_15_output_z_ack;

	wire [31:0] adder_15_output_z;
	wire adder_15_output_z_stb;
	wire adder_15_input_a_ack;
	wire adder_15_input_b_ack;

	reg	[1:0] adder_15_state;
parameter adder_15_put_a         = 2'd0,
          adder_15_put_b         = 2'd1,
          adder_15_get_z         = 2'd2;
	adder_15 adder_15_inst (adder_15_input_a, adder_15_input_b, adder_15_input_a_stb, adder_15_input_b_stb, adder_15_output_z_ack, clock_signal, reset_signal, adder_15_output_z, adder_15_output_z_stb, adder_15_input_a_ack, adder_15_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_15_input_a;
	reg [31:0] multiplier_15_input_b;
	reg multiplier_15_input_a_stb;
	reg multiplier_15_input_b_stb;
	reg multiplier_15_output_z_ack;

	wire [31:0] multiplier_15_output_z;
	wire multiplier_15_output_z_stb;
	wire multiplier_15_input_a_ack;
	wire multiplier_15_input_b_ack;

	reg	[1:0] multiplier_15_state;
parameter multiplier_15_put_a         = 2'd0,
          multiplier_15_put_b         = 2'd1,
          multiplier_15_get_z         = 2'd2;
	multiplier_15 multiplier_15_inst (multiplier_15_input_a, multiplier_15_input_b, multiplier_15_input_a_stb, multiplier_15_input_b_stb, multiplier_15_output_z_ack, clock_signal, reset_signal, multiplier_15_output_z, multiplier_15_output_z_stb, multiplier_15_input_a_ack, multiplier_15_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_15_state)
							adder_15_put_a : begin
								if (adder_15_input_a_ack) begin
									adder_15_input_a <= #1 _r0;
									adder_15_input_a_stb <= #1 1;
									adder_15_output_z_ack <= #1 0;
									adder_15_state <= #1 adder_15_put_b;
								end
							end
							adder_15_put_b : begin
								if (adder_15_input_b_ack) begin
									adder_15_input_b <= #1 _r7;
									adder_15_input_b_stb <= #1 1;
									adder_15_output_z_ack <= #1 0;
									adder_15_state <= #1 adder_15_get_z;
									adder_15_input_a_stb <= #1 0;
								end
							end
							adder_15_get_z : begin
								if (adder_15_output_z_stb) begin
									_r0 <= #1 adder_15_output_z;
									adder_15_output_z_ack <= #1 1;
									adder_15_state <= #1 adder_15_put_a;
									adder_15_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_15_state)
							adder_15_put_a : begin
								if (adder_15_input_a_ack) begin
									adder_15_input_a <= #1 _r6;
									adder_15_input_a_stb <= #1 1;
									adder_15_output_z_ack <= #1 0;
									adder_15_state <= #1 adder_15_put_b;
								end
							end
							adder_15_put_b : begin
								if (adder_15_input_b_ack) begin
									adder_15_input_b <= #1 _r7;
									adder_15_input_b_stb <= #1 1;
									adder_15_output_z_ack <= #1 0;
									adder_15_state <= #1 adder_15_get_z;
									adder_15_input_a_stb <= #1 0;
								end
							end
							adder_15_get_z : begin
								if (adder_15_output_z_stb) begin
									_r6 <= #1 adder_15_output_z;
									adder_15_output_z_ack <= #1 1;
									adder_15_state <= #1 adder_15_put_a;
									adder_15_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_15_state)
							multiplier_15_put_a : begin
								if (multiplier_15_input_a_ack) begin
									multiplier_15_input_a <= #1 _r0;
									multiplier_15_input_a_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_put_b;
								end
							end
							multiplier_15_put_b : begin
								if (multiplier_15_input_b_ack) begin
									multiplier_15_input_b <= #1 _r3;
									multiplier_15_input_b_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_get_z;
									multiplier_15_input_a_stb <= #1 0;
								end
							end
							multiplier_15_get_z : begin
								if (multiplier_15_output_z_stb) begin
									_r0 <= #1 multiplier_15_output_z;
									multiplier_15_output_z_ack <= #1 1;
									multiplier_15_state <= #1 multiplier_15_put_a;
									multiplier_15_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_15_state)
							multiplier_15_put_a : begin
								if (multiplier_15_input_a_ack) begin
									multiplier_15_input_a <= #1 _r0;
									multiplier_15_input_a_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_put_b;
								end
							end
							multiplier_15_put_b : begin
								if (multiplier_15_input_b_ack) begin
									multiplier_15_input_b <= #1 _r4;
									multiplier_15_input_b_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_get_z;
									multiplier_15_input_a_stb <= #1 0;
								end
							end
							multiplier_15_get_z : begin
								if (multiplier_15_output_z_stb) begin
									_r0 <= #1 multiplier_15_output_z;
									multiplier_15_output_z_ack <= #1 1;
									multiplier_15_state <= #1 multiplier_15_put_a;
									multiplier_15_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_15_state)
							multiplier_15_put_a : begin
								if (multiplier_15_input_a_ack) begin
									multiplier_15_input_a <= #1 _r0;
									multiplier_15_input_a_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_put_b;
								end
							end
							multiplier_15_put_b : begin
								if (multiplier_15_input_b_ack) begin
									multiplier_15_input_b <= #1 _r5;
									multiplier_15_input_b_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_get_z;
									multiplier_15_input_a_stb <= #1 0;
								end
							end
							multiplier_15_get_z : begin
								if (multiplier_15_output_z_stb) begin
									_r0 <= #1 multiplier_15_output_z;
									multiplier_15_output_z_ack <= #1 1;
									multiplier_15_state <= #1 multiplier_15_put_a;
									multiplier_15_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_15_state)
							multiplier_15_put_a : begin
								if (multiplier_15_input_a_ack) begin
									multiplier_15_input_a <= #1 _r7;
									multiplier_15_input_a_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_put_b;
								end
							end
							multiplier_15_put_b : begin
								if (multiplier_15_input_b_ack) begin
									multiplier_15_input_b <= #1 _r3;
									multiplier_15_input_b_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_get_z;
									multiplier_15_input_a_stb <= #1 0;
								end
							end
							multiplier_15_get_z : begin
								if (multiplier_15_output_z_stb) begin
									_r7 <= #1 multiplier_15_output_z;
									multiplier_15_output_z_ack <= #1 1;
									multiplier_15_state <= #1 multiplier_15_put_a;
									multiplier_15_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_15_state)
							multiplier_15_put_a : begin
								if (multiplier_15_input_a_ack) begin
									multiplier_15_input_a <= #1 _r7;
									multiplier_15_input_a_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_put_b;
								end
							end
							multiplier_15_put_b : begin
								if (multiplier_15_input_b_ack) begin
									multiplier_15_input_b <= #1 _r4;
									multiplier_15_input_b_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_get_z;
									multiplier_15_input_a_stb <= #1 0;
								end
							end
							multiplier_15_get_z : begin
								if (multiplier_15_output_z_stb) begin
									_r7 <= #1 multiplier_15_output_z;
									multiplier_15_output_z_ack <= #1 1;
									multiplier_15_state <= #1 multiplier_15_put_a;
									multiplier_15_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_15_state)
							multiplier_15_put_a : begin
								if (multiplier_15_input_a_ack) begin
									multiplier_15_input_a <= #1 _r7;
									multiplier_15_input_a_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_put_b;
								end
							end
							multiplier_15_put_b : begin
								if (multiplier_15_input_b_ack) begin
									multiplier_15_input_b <= #1 _r5;
									multiplier_15_input_b_stb <= #1 1;
									multiplier_15_output_z_ack <= #1 0;
									multiplier_15_state <= #1 multiplier_15_get_z;
									multiplier_15_input_a_stb <= #1 0;
								end
							end
							multiplier_15_get_z : begin
								if (multiplier_15_output_z_stb) begin
									_r7 <= #1 multiplier_15_output_z;
									multiplier_15_output_z_ack <= #1 1;
									multiplier_15_state <= #1 multiplier_15_put_a;
									multiplier_15_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_15 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_15 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p16ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b10000000000000000000000000000000;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00111111100000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p16rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p16(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_16_input_a;
	reg [31:0] adder_16_input_b;
	reg adder_16_input_a_stb;
	reg adder_16_input_b_stb;
	reg adder_16_output_z_ack;

	wire [31:0] adder_16_output_z;
	wire adder_16_output_z_stb;
	wire adder_16_input_a_ack;
	wire adder_16_input_b_ack;

	reg	[1:0] adder_16_state;
parameter adder_16_put_a         = 2'd0,
          adder_16_put_b         = 2'd1,
          adder_16_get_z         = 2'd2;
	adder_16 adder_16_inst (adder_16_input_a, adder_16_input_b, adder_16_input_a_stb, adder_16_input_b_stb, adder_16_output_z_ack, clock_signal, reset_signal, adder_16_output_z, adder_16_output_z_stb, adder_16_input_a_ack, adder_16_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_16_input_a;
	reg [31:0] multiplier_16_input_b;
	reg multiplier_16_input_a_stb;
	reg multiplier_16_input_b_stb;
	reg multiplier_16_output_z_ack;

	wire [31:0] multiplier_16_output_z;
	wire multiplier_16_output_z_stb;
	wire multiplier_16_input_a_ack;
	wire multiplier_16_input_b_ack;

	reg	[1:0] multiplier_16_state;
parameter multiplier_16_put_a         = 2'd0,
          multiplier_16_put_b         = 2'd1,
          multiplier_16_get_z         = 2'd2;
	multiplier_16 multiplier_16_inst (multiplier_16_input_a, multiplier_16_input_b, multiplier_16_input_a_stb, multiplier_16_input_b_stb, multiplier_16_output_z_ack, clock_signal, reset_signal, multiplier_16_output_z, multiplier_16_output_z_stb, multiplier_16_input_a_ack, multiplier_16_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_16_state)
							adder_16_put_a : begin
								if (adder_16_input_a_ack) begin
									adder_16_input_a <= #1 _r0;
									adder_16_input_a_stb <= #1 1;
									adder_16_output_z_ack <= #1 0;
									adder_16_state <= #1 adder_16_put_b;
								end
							end
							adder_16_put_b : begin
								if (adder_16_input_b_ack) begin
									adder_16_input_b <= #1 _r7;
									adder_16_input_b_stb <= #1 1;
									adder_16_output_z_ack <= #1 0;
									adder_16_state <= #1 adder_16_get_z;
									adder_16_input_a_stb <= #1 0;
								end
							end
							adder_16_get_z : begin
								if (adder_16_output_z_stb) begin
									_r0 <= #1 adder_16_output_z;
									adder_16_output_z_ack <= #1 1;
									adder_16_state <= #1 adder_16_put_a;
									adder_16_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_16_state)
							adder_16_put_a : begin
								if (adder_16_input_a_ack) begin
									adder_16_input_a <= #1 _r6;
									adder_16_input_a_stb <= #1 1;
									adder_16_output_z_ack <= #1 0;
									adder_16_state <= #1 adder_16_put_b;
								end
							end
							adder_16_put_b : begin
								if (adder_16_input_b_ack) begin
									adder_16_input_b <= #1 _r7;
									adder_16_input_b_stb <= #1 1;
									adder_16_output_z_ack <= #1 0;
									adder_16_state <= #1 adder_16_get_z;
									adder_16_input_a_stb <= #1 0;
								end
							end
							adder_16_get_z : begin
								if (adder_16_output_z_stb) begin
									_r6 <= #1 adder_16_output_z;
									adder_16_output_z_ack <= #1 1;
									adder_16_state <= #1 adder_16_put_a;
									adder_16_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_16_state)
							multiplier_16_put_a : begin
								if (multiplier_16_input_a_ack) begin
									multiplier_16_input_a <= #1 _r0;
									multiplier_16_input_a_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_put_b;
								end
							end
							multiplier_16_put_b : begin
								if (multiplier_16_input_b_ack) begin
									multiplier_16_input_b <= #1 _r3;
									multiplier_16_input_b_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_get_z;
									multiplier_16_input_a_stb <= #1 0;
								end
							end
							multiplier_16_get_z : begin
								if (multiplier_16_output_z_stb) begin
									_r0 <= #1 multiplier_16_output_z;
									multiplier_16_output_z_ack <= #1 1;
									multiplier_16_state <= #1 multiplier_16_put_a;
									multiplier_16_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_16_state)
							multiplier_16_put_a : begin
								if (multiplier_16_input_a_ack) begin
									multiplier_16_input_a <= #1 _r0;
									multiplier_16_input_a_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_put_b;
								end
							end
							multiplier_16_put_b : begin
								if (multiplier_16_input_b_ack) begin
									multiplier_16_input_b <= #1 _r4;
									multiplier_16_input_b_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_get_z;
									multiplier_16_input_a_stb <= #1 0;
								end
							end
							multiplier_16_get_z : begin
								if (multiplier_16_output_z_stb) begin
									_r0 <= #1 multiplier_16_output_z;
									multiplier_16_output_z_ack <= #1 1;
									multiplier_16_state <= #1 multiplier_16_put_a;
									multiplier_16_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_16_state)
							multiplier_16_put_a : begin
								if (multiplier_16_input_a_ack) begin
									multiplier_16_input_a <= #1 _r0;
									multiplier_16_input_a_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_put_b;
								end
							end
							multiplier_16_put_b : begin
								if (multiplier_16_input_b_ack) begin
									multiplier_16_input_b <= #1 _r5;
									multiplier_16_input_b_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_get_z;
									multiplier_16_input_a_stb <= #1 0;
								end
							end
							multiplier_16_get_z : begin
								if (multiplier_16_output_z_stb) begin
									_r0 <= #1 multiplier_16_output_z;
									multiplier_16_output_z_ack <= #1 1;
									multiplier_16_state <= #1 multiplier_16_put_a;
									multiplier_16_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_16_state)
							multiplier_16_put_a : begin
								if (multiplier_16_input_a_ack) begin
									multiplier_16_input_a <= #1 _r7;
									multiplier_16_input_a_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_put_b;
								end
							end
							multiplier_16_put_b : begin
								if (multiplier_16_input_b_ack) begin
									multiplier_16_input_b <= #1 _r3;
									multiplier_16_input_b_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_get_z;
									multiplier_16_input_a_stb <= #1 0;
								end
							end
							multiplier_16_get_z : begin
								if (multiplier_16_output_z_stb) begin
									_r7 <= #1 multiplier_16_output_z;
									multiplier_16_output_z_ack <= #1 1;
									multiplier_16_state <= #1 multiplier_16_put_a;
									multiplier_16_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_16_state)
							multiplier_16_put_a : begin
								if (multiplier_16_input_a_ack) begin
									multiplier_16_input_a <= #1 _r7;
									multiplier_16_input_a_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_put_b;
								end
							end
							multiplier_16_put_b : begin
								if (multiplier_16_input_b_ack) begin
									multiplier_16_input_b <= #1 _r4;
									multiplier_16_input_b_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_get_z;
									multiplier_16_input_a_stb <= #1 0;
								end
							end
							multiplier_16_get_z : begin
								if (multiplier_16_output_z_stb) begin
									_r7 <= #1 multiplier_16_output_z;
									multiplier_16_output_z_ack <= #1 1;
									multiplier_16_state <= #1 multiplier_16_put_a;
									multiplier_16_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_16_state)
							multiplier_16_put_a : begin
								if (multiplier_16_input_a_ack) begin
									multiplier_16_input_a <= #1 _r7;
									multiplier_16_input_a_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_put_b;
								end
							end
							multiplier_16_put_b : begin
								if (multiplier_16_input_b_ack) begin
									multiplier_16_input_b <= #1 _r5;
									multiplier_16_input_b_stb <= #1 1;
									multiplier_16_output_z_ack <= #1 0;
									multiplier_16_state <= #1 multiplier_16_get_z;
									multiplier_16_input_a_stb <= #1 0;
								end
							end
							multiplier_16_get_z : begin
								if (multiplier_16_output_z_stb) begin
									_r7 <= #1 multiplier_16_output_z;
									multiplier_16_output_z_ack <= #1 1;
									multiplier_16_state <= #1 multiplier_16_put_a;
									multiplier_16_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_16 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_16 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p17ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00000000000000000000000000000000;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p17rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p17(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_17_input_a;
	reg [31:0] adder_17_input_b;
	reg adder_17_input_a_stb;
	reg adder_17_input_b_stb;
	reg adder_17_output_z_ack;

	wire [31:0] adder_17_output_z;
	wire adder_17_output_z_stb;
	wire adder_17_input_a_ack;
	wire adder_17_input_b_ack;

	reg	[1:0] adder_17_state;
parameter adder_17_put_a         = 2'd0,
          adder_17_put_b         = 2'd1,
          adder_17_get_z         = 2'd2;
	adder_17 adder_17_inst (adder_17_input_a, adder_17_input_b, adder_17_input_a_stb, adder_17_input_b_stb, adder_17_output_z_ack, clock_signal, reset_signal, adder_17_output_z, adder_17_output_z_stb, adder_17_input_a_ack, adder_17_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_17_input_a;
	reg [31:0] multiplier_17_input_b;
	reg multiplier_17_input_a_stb;
	reg multiplier_17_input_b_stb;
	reg multiplier_17_output_z_ack;

	wire [31:0] multiplier_17_output_z;
	wire multiplier_17_output_z_stb;
	wire multiplier_17_input_a_ack;
	wire multiplier_17_input_b_ack;

	reg	[1:0] multiplier_17_state;
parameter multiplier_17_put_a         = 2'd0,
          multiplier_17_put_b         = 2'd1,
          multiplier_17_get_z         = 2'd2;
	multiplier_17 multiplier_17_inst (multiplier_17_input_a, multiplier_17_input_b, multiplier_17_input_a_stb, multiplier_17_input_b_stb, multiplier_17_output_z_ack, clock_signal, reset_signal, multiplier_17_output_z, multiplier_17_output_z_stb, multiplier_17_input_a_ack, multiplier_17_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_17_state)
							adder_17_put_a : begin
								if (adder_17_input_a_ack) begin
									adder_17_input_a <= #1 _r0;
									adder_17_input_a_stb <= #1 1;
									adder_17_output_z_ack <= #1 0;
									adder_17_state <= #1 adder_17_put_b;
								end
							end
							adder_17_put_b : begin
								if (adder_17_input_b_ack) begin
									adder_17_input_b <= #1 _r7;
									adder_17_input_b_stb <= #1 1;
									adder_17_output_z_ack <= #1 0;
									adder_17_state <= #1 adder_17_get_z;
									adder_17_input_a_stb <= #1 0;
								end
							end
							adder_17_get_z : begin
								if (adder_17_output_z_stb) begin
									_r0 <= #1 adder_17_output_z;
									adder_17_output_z_ack <= #1 1;
									adder_17_state <= #1 adder_17_put_a;
									adder_17_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_17_state)
							adder_17_put_a : begin
								if (adder_17_input_a_ack) begin
									adder_17_input_a <= #1 _r6;
									adder_17_input_a_stb <= #1 1;
									adder_17_output_z_ack <= #1 0;
									adder_17_state <= #1 adder_17_put_b;
								end
							end
							adder_17_put_b : begin
								if (adder_17_input_b_ack) begin
									adder_17_input_b <= #1 _r7;
									adder_17_input_b_stb <= #1 1;
									adder_17_output_z_ack <= #1 0;
									adder_17_state <= #1 adder_17_get_z;
									adder_17_input_a_stb <= #1 0;
								end
							end
							adder_17_get_z : begin
								if (adder_17_output_z_stb) begin
									_r6 <= #1 adder_17_output_z;
									adder_17_output_z_ack <= #1 1;
									adder_17_state <= #1 adder_17_put_a;
									adder_17_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_17_state)
							multiplier_17_put_a : begin
								if (multiplier_17_input_a_ack) begin
									multiplier_17_input_a <= #1 _r0;
									multiplier_17_input_a_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_put_b;
								end
							end
							multiplier_17_put_b : begin
								if (multiplier_17_input_b_ack) begin
									multiplier_17_input_b <= #1 _r3;
									multiplier_17_input_b_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_get_z;
									multiplier_17_input_a_stb <= #1 0;
								end
							end
							multiplier_17_get_z : begin
								if (multiplier_17_output_z_stb) begin
									_r0 <= #1 multiplier_17_output_z;
									multiplier_17_output_z_ack <= #1 1;
									multiplier_17_state <= #1 multiplier_17_put_a;
									multiplier_17_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_17_state)
							multiplier_17_put_a : begin
								if (multiplier_17_input_a_ack) begin
									multiplier_17_input_a <= #1 _r0;
									multiplier_17_input_a_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_put_b;
								end
							end
							multiplier_17_put_b : begin
								if (multiplier_17_input_b_ack) begin
									multiplier_17_input_b <= #1 _r4;
									multiplier_17_input_b_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_get_z;
									multiplier_17_input_a_stb <= #1 0;
								end
							end
							multiplier_17_get_z : begin
								if (multiplier_17_output_z_stb) begin
									_r0 <= #1 multiplier_17_output_z;
									multiplier_17_output_z_ack <= #1 1;
									multiplier_17_state <= #1 multiplier_17_put_a;
									multiplier_17_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_17_state)
							multiplier_17_put_a : begin
								if (multiplier_17_input_a_ack) begin
									multiplier_17_input_a <= #1 _r0;
									multiplier_17_input_a_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_put_b;
								end
							end
							multiplier_17_put_b : begin
								if (multiplier_17_input_b_ack) begin
									multiplier_17_input_b <= #1 _r5;
									multiplier_17_input_b_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_get_z;
									multiplier_17_input_a_stb <= #1 0;
								end
							end
							multiplier_17_get_z : begin
								if (multiplier_17_output_z_stb) begin
									_r0 <= #1 multiplier_17_output_z;
									multiplier_17_output_z_ack <= #1 1;
									multiplier_17_state <= #1 multiplier_17_put_a;
									multiplier_17_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_17_state)
							multiplier_17_put_a : begin
								if (multiplier_17_input_a_ack) begin
									multiplier_17_input_a <= #1 _r7;
									multiplier_17_input_a_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_put_b;
								end
							end
							multiplier_17_put_b : begin
								if (multiplier_17_input_b_ack) begin
									multiplier_17_input_b <= #1 _r3;
									multiplier_17_input_b_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_get_z;
									multiplier_17_input_a_stb <= #1 0;
								end
							end
							multiplier_17_get_z : begin
								if (multiplier_17_output_z_stb) begin
									_r7 <= #1 multiplier_17_output_z;
									multiplier_17_output_z_ack <= #1 1;
									multiplier_17_state <= #1 multiplier_17_put_a;
									multiplier_17_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_17_state)
							multiplier_17_put_a : begin
								if (multiplier_17_input_a_ack) begin
									multiplier_17_input_a <= #1 _r7;
									multiplier_17_input_a_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_put_b;
								end
							end
							multiplier_17_put_b : begin
								if (multiplier_17_input_b_ack) begin
									multiplier_17_input_b <= #1 _r4;
									multiplier_17_input_b_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_get_z;
									multiplier_17_input_a_stb <= #1 0;
								end
							end
							multiplier_17_get_z : begin
								if (multiplier_17_output_z_stb) begin
									_r7 <= #1 multiplier_17_output_z;
									multiplier_17_output_z_ack <= #1 1;
									multiplier_17_state <= #1 multiplier_17_put_a;
									multiplier_17_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_17_state)
							multiplier_17_put_a : begin
								if (multiplier_17_input_a_ack) begin
									multiplier_17_input_a <= #1 _r7;
									multiplier_17_input_a_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_put_b;
								end
							end
							multiplier_17_put_b : begin
								if (multiplier_17_input_b_ack) begin
									multiplier_17_input_b <= #1 _r5;
									multiplier_17_input_b_stb <= #1 1;
									multiplier_17_output_z_ack <= #1 0;
									multiplier_17_state <= #1 multiplier_17_get_z;
									multiplier_17_input_a_stb <= #1 0;
								end
							end
							multiplier_17_get_z : begin
								if (multiplier_17_output_z_stb) begin
									_r7 <= #1 multiplier_17_output_z;
									multiplier_17_output_z_ack <= #1 1;
									multiplier_17_state <= #1 multiplier_17_put_a;
									multiplier_17_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_17 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_17 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p18ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00111111001101010000010011110011;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p18rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p18(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_18_input_a;
	reg [31:0] adder_18_input_b;
	reg adder_18_input_a_stb;
	reg adder_18_input_b_stb;
	reg adder_18_output_z_ack;

	wire [31:0] adder_18_output_z;
	wire adder_18_output_z_stb;
	wire adder_18_input_a_ack;
	wire adder_18_input_b_ack;

	reg	[1:0] adder_18_state;
parameter adder_18_put_a         = 2'd0,
          adder_18_put_b         = 2'd1,
          adder_18_get_z         = 2'd2;
	adder_18 adder_18_inst (adder_18_input_a, adder_18_input_b, adder_18_input_a_stb, adder_18_input_b_stb, adder_18_output_z_ack, clock_signal, reset_signal, adder_18_output_z, adder_18_output_z_stb, adder_18_input_a_ack, adder_18_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_18_input_a;
	reg [31:0] multiplier_18_input_b;
	reg multiplier_18_input_a_stb;
	reg multiplier_18_input_b_stb;
	reg multiplier_18_output_z_ack;

	wire [31:0] multiplier_18_output_z;
	wire multiplier_18_output_z_stb;
	wire multiplier_18_input_a_ack;
	wire multiplier_18_input_b_ack;

	reg	[1:0] multiplier_18_state;
parameter multiplier_18_put_a         = 2'd0,
          multiplier_18_put_b         = 2'd1,
          multiplier_18_get_z         = 2'd2;
	multiplier_18 multiplier_18_inst (multiplier_18_input_a, multiplier_18_input_b, multiplier_18_input_a_stb, multiplier_18_input_b_stb, multiplier_18_output_z_ack, clock_signal, reset_signal, multiplier_18_output_z, multiplier_18_output_z_stb, multiplier_18_input_a_ack, multiplier_18_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_18_state)
							adder_18_put_a : begin
								if (adder_18_input_a_ack) begin
									adder_18_input_a <= #1 _r0;
									adder_18_input_a_stb <= #1 1;
									adder_18_output_z_ack <= #1 0;
									adder_18_state <= #1 adder_18_put_b;
								end
							end
							adder_18_put_b : begin
								if (adder_18_input_b_ack) begin
									adder_18_input_b <= #1 _r7;
									adder_18_input_b_stb <= #1 1;
									adder_18_output_z_ack <= #1 0;
									adder_18_state <= #1 adder_18_get_z;
									adder_18_input_a_stb <= #1 0;
								end
							end
							adder_18_get_z : begin
								if (adder_18_output_z_stb) begin
									_r0 <= #1 adder_18_output_z;
									adder_18_output_z_ack <= #1 1;
									adder_18_state <= #1 adder_18_put_a;
									adder_18_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_18_state)
							adder_18_put_a : begin
								if (adder_18_input_a_ack) begin
									adder_18_input_a <= #1 _r6;
									adder_18_input_a_stb <= #1 1;
									adder_18_output_z_ack <= #1 0;
									adder_18_state <= #1 adder_18_put_b;
								end
							end
							adder_18_put_b : begin
								if (adder_18_input_b_ack) begin
									adder_18_input_b <= #1 _r7;
									adder_18_input_b_stb <= #1 1;
									adder_18_output_z_ack <= #1 0;
									adder_18_state <= #1 adder_18_get_z;
									adder_18_input_a_stb <= #1 0;
								end
							end
							adder_18_get_z : begin
								if (adder_18_output_z_stb) begin
									_r6 <= #1 adder_18_output_z;
									adder_18_output_z_ack <= #1 1;
									adder_18_state <= #1 adder_18_put_a;
									adder_18_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_18_state)
							multiplier_18_put_a : begin
								if (multiplier_18_input_a_ack) begin
									multiplier_18_input_a <= #1 _r0;
									multiplier_18_input_a_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_put_b;
								end
							end
							multiplier_18_put_b : begin
								if (multiplier_18_input_b_ack) begin
									multiplier_18_input_b <= #1 _r3;
									multiplier_18_input_b_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_get_z;
									multiplier_18_input_a_stb <= #1 0;
								end
							end
							multiplier_18_get_z : begin
								if (multiplier_18_output_z_stb) begin
									_r0 <= #1 multiplier_18_output_z;
									multiplier_18_output_z_ack <= #1 1;
									multiplier_18_state <= #1 multiplier_18_put_a;
									multiplier_18_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_18_state)
							multiplier_18_put_a : begin
								if (multiplier_18_input_a_ack) begin
									multiplier_18_input_a <= #1 _r0;
									multiplier_18_input_a_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_put_b;
								end
							end
							multiplier_18_put_b : begin
								if (multiplier_18_input_b_ack) begin
									multiplier_18_input_b <= #1 _r4;
									multiplier_18_input_b_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_get_z;
									multiplier_18_input_a_stb <= #1 0;
								end
							end
							multiplier_18_get_z : begin
								if (multiplier_18_output_z_stb) begin
									_r0 <= #1 multiplier_18_output_z;
									multiplier_18_output_z_ack <= #1 1;
									multiplier_18_state <= #1 multiplier_18_put_a;
									multiplier_18_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_18_state)
							multiplier_18_put_a : begin
								if (multiplier_18_input_a_ack) begin
									multiplier_18_input_a <= #1 _r0;
									multiplier_18_input_a_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_put_b;
								end
							end
							multiplier_18_put_b : begin
								if (multiplier_18_input_b_ack) begin
									multiplier_18_input_b <= #1 _r5;
									multiplier_18_input_b_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_get_z;
									multiplier_18_input_a_stb <= #1 0;
								end
							end
							multiplier_18_get_z : begin
								if (multiplier_18_output_z_stb) begin
									_r0 <= #1 multiplier_18_output_z;
									multiplier_18_output_z_ack <= #1 1;
									multiplier_18_state <= #1 multiplier_18_put_a;
									multiplier_18_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_18_state)
							multiplier_18_put_a : begin
								if (multiplier_18_input_a_ack) begin
									multiplier_18_input_a <= #1 _r7;
									multiplier_18_input_a_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_put_b;
								end
							end
							multiplier_18_put_b : begin
								if (multiplier_18_input_b_ack) begin
									multiplier_18_input_b <= #1 _r3;
									multiplier_18_input_b_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_get_z;
									multiplier_18_input_a_stb <= #1 0;
								end
							end
							multiplier_18_get_z : begin
								if (multiplier_18_output_z_stb) begin
									_r7 <= #1 multiplier_18_output_z;
									multiplier_18_output_z_ack <= #1 1;
									multiplier_18_state <= #1 multiplier_18_put_a;
									multiplier_18_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_18_state)
							multiplier_18_put_a : begin
								if (multiplier_18_input_a_ack) begin
									multiplier_18_input_a <= #1 _r7;
									multiplier_18_input_a_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_put_b;
								end
							end
							multiplier_18_put_b : begin
								if (multiplier_18_input_b_ack) begin
									multiplier_18_input_b <= #1 _r4;
									multiplier_18_input_b_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_get_z;
									multiplier_18_input_a_stb <= #1 0;
								end
							end
							multiplier_18_get_z : begin
								if (multiplier_18_output_z_stb) begin
									_r7 <= #1 multiplier_18_output_z;
									multiplier_18_output_z_ack <= #1 1;
									multiplier_18_state <= #1 multiplier_18_put_a;
									multiplier_18_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_18_state)
							multiplier_18_put_a : begin
								if (multiplier_18_input_a_ack) begin
									multiplier_18_input_a <= #1 _r7;
									multiplier_18_input_a_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_put_b;
								end
							end
							multiplier_18_put_b : begin
								if (multiplier_18_input_b_ack) begin
									multiplier_18_input_b <= #1 _r5;
									multiplier_18_input_b_stb <= #1 1;
									multiplier_18_output_z_ack <= #1 0;
									multiplier_18_state <= #1 multiplier_18_get_z;
									multiplier_18_input_a_stb <= #1 0;
								end
							end
							multiplier_18_get_z : begin
								if (multiplier_18_output_z_stb) begin
									_r7 <= #1 multiplier_18_output_z;
									multiplier_18_output_z_ack <= #1 1;
									multiplier_18_state <= #1 multiplier_18_put_a;
									multiplier_18_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_18 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_18 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p19ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b10000000000000000000000000000000;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00111111100000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p19rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p19(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_19_input_a;
	reg [31:0] adder_19_input_b;
	reg adder_19_input_a_stb;
	reg adder_19_input_b_stb;
	reg adder_19_output_z_ack;

	wire [31:0] adder_19_output_z;
	wire adder_19_output_z_stb;
	wire adder_19_input_a_ack;
	wire adder_19_input_b_ack;

	reg	[1:0] adder_19_state;
parameter adder_19_put_a         = 2'd0,
          adder_19_put_b         = 2'd1,
          adder_19_get_z         = 2'd2;
	adder_19 adder_19_inst (adder_19_input_a, adder_19_input_b, adder_19_input_a_stb, adder_19_input_b_stb, adder_19_output_z_ack, clock_signal, reset_signal, adder_19_output_z, adder_19_output_z_stb, adder_19_input_a_ack, adder_19_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_19_input_a;
	reg [31:0] multiplier_19_input_b;
	reg multiplier_19_input_a_stb;
	reg multiplier_19_input_b_stb;
	reg multiplier_19_output_z_ack;

	wire [31:0] multiplier_19_output_z;
	wire multiplier_19_output_z_stb;
	wire multiplier_19_input_a_ack;
	wire multiplier_19_input_b_ack;

	reg	[1:0] multiplier_19_state;
parameter multiplier_19_put_a         = 2'd0,
          multiplier_19_put_b         = 2'd1,
          multiplier_19_get_z         = 2'd2;
	multiplier_19 multiplier_19_inst (multiplier_19_input_a, multiplier_19_input_b, multiplier_19_input_a_stb, multiplier_19_input_b_stb, multiplier_19_output_z_ack, clock_signal, reset_signal, multiplier_19_output_z, multiplier_19_output_z_stb, multiplier_19_input_a_ack, multiplier_19_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_19_state)
							adder_19_put_a : begin
								if (adder_19_input_a_ack) begin
									adder_19_input_a <= #1 _r0;
									adder_19_input_a_stb <= #1 1;
									adder_19_output_z_ack <= #1 0;
									adder_19_state <= #1 adder_19_put_b;
								end
							end
							adder_19_put_b : begin
								if (adder_19_input_b_ack) begin
									adder_19_input_b <= #1 _r7;
									adder_19_input_b_stb <= #1 1;
									adder_19_output_z_ack <= #1 0;
									adder_19_state <= #1 adder_19_get_z;
									adder_19_input_a_stb <= #1 0;
								end
							end
							adder_19_get_z : begin
								if (adder_19_output_z_stb) begin
									_r0 <= #1 adder_19_output_z;
									adder_19_output_z_ack <= #1 1;
									adder_19_state <= #1 adder_19_put_a;
									adder_19_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_19_state)
							adder_19_put_a : begin
								if (adder_19_input_a_ack) begin
									adder_19_input_a <= #1 _r6;
									adder_19_input_a_stb <= #1 1;
									adder_19_output_z_ack <= #1 0;
									adder_19_state <= #1 adder_19_put_b;
								end
							end
							adder_19_put_b : begin
								if (adder_19_input_b_ack) begin
									adder_19_input_b <= #1 _r7;
									adder_19_input_b_stb <= #1 1;
									adder_19_output_z_ack <= #1 0;
									adder_19_state <= #1 adder_19_get_z;
									adder_19_input_a_stb <= #1 0;
								end
							end
							adder_19_get_z : begin
								if (adder_19_output_z_stb) begin
									_r6 <= #1 adder_19_output_z;
									adder_19_output_z_ack <= #1 1;
									adder_19_state <= #1 adder_19_put_a;
									adder_19_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_19_state)
							multiplier_19_put_a : begin
								if (multiplier_19_input_a_ack) begin
									multiplier_19_input_a <= #1 _r0;
									multiplier_19_input_a_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_put_b;
								end
							end
							multiplier_19_put_b : begin
								if (multiplier_19_input_b_ack) begin
									multiplier_19_input_b <= #1 _r3;
									multiplier_19_input_b_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_get_z;
									multiplier_19_input_a_stb <= #1 0;
								end
							end
							multiplier_19_get_z : begin
								if (multiplier_19_output_z_stb) begin
									_r0 <= #1 multiplier_19_output_z;
									multiplier_19_output_z_ack <= #1 1;
									multiplier_19_state <= #1 multiplier_19_put_a;
									multiplier_19_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_19_state)
							multiplier_19_put_a : begin
								if (multiplier_19_input_a_ack) begin
									multiplier_19_input_a <= #1 _r0;
									multiplier_19_input_a_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_put_b;
								end
							end
							multiplier_19_put_b : begin
								if (multiplier_19_input_b_ack) begin
									multiplier_19_input_b <= #1 _r4;
									multiplier_19_input_b_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_get_z;
									multiplier_19_input_a_stb <= #1 0;
								end
							end
							multiplier_19_get_z : begin
								if (multiplier_19_output_z_stb) begin
									_r0 <= #1 multiplier_19_output_z;
									multiplier_19_output_z_ack <= #1 1;
									multiplier_19_state <= #1 multiplier_19_put_a;
									multiplier_19_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_19_state)
							multiplier_19_put_a : begin
								if (multiplier_19_input_a_ack) begin
									multiplier_19_input_a <= #1 _r0;
									multiplier_19_input_a_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_put_b;
								end
							end
							multiplier_19_put_b : begin
								if (multiplier_19_input_b_ack) begin
									multiplier_19_input_b <= #1 _r5;
									multiplier_19_input_b_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_get_z;
									multiplier_19_input_a_stb <= #1 0;
								end
							end
							multiplier_19_get_z : begin
								if (multiplier_19_output_z_stb) begin
									_r0 <= #1 multiplier_19_output_z;
									multiplier_19_output_z_ack <= #1 1;
									multiplier_19_state <= #1 multiplier_19_put_a;
									multiplier_19_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_19_state)
							multiplier_19_put_a : begin
								if (multiplier_19_input_a_ack) begin
									multiplier_19_input_a <= #1 _r7;
									multiplier_19_input_a_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_put_b;
								end
							end
							multiplier_19_put_b : begin
								if (multiplier_19_input_b_ack) begin
									multiplier_19_input_b <= #1 _r3;
									multiplier_19_input_b_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_get_z;
									multiplier_19_input_a_stb <= #1 0;
								end
							end
							multiplier_19_get_z : begin
								if (multiplier_19_output_z_stb) begin
									_r7 <= #1 multiplier_19_output_z;
									multiplier_19_output_z_ack <= #1 1;
									multiplier_19_state <= #1 multiplier_19_put_a;
									multiplier_19_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_19_state)
							multiplier_19_put_a : begin
								if (multiplier_19_input_a_ack) begin
									multiplier_19_input_a <= #1 _r7;
									multiplier_19_input_a_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_put_b;
								end
							end
							multiplier_19_put_b : begin
								if (multiplier_19_input_b_ack) begin
									multiplier_19_input_b <= #1 _r4;
									multiplier_19_input_b_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_get_z;
									multiplier_19_input_a_stb <= #1 0;
								end
							end
							multiplier_19_get_z : begin
								if (multiplier_19_output_z_stb) begin
									_r7 <= #1 multiplier_19_output_z;
									multiplier_19_output_z_ack <= #1 1;
									multiplier_19_state <= #1 multiplier_19_put_a;
									multiplier_19_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_19_state)
							multiplier_19_put_a : begin
								if (multiplier_19_input_a_ack) begin
									multiplier_19_input_a <= #1 _r7;
									multiplier_19_input_a_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_put_b;
								end
							end
							multiplier_19_put_b : begin
								if (multiplier_19_input_b_ack) begin
									multiplier_19_input_b <= #1 _r5;
									multiplier_19_input_b_stb <= #1 1;
									multiplier_19_output_z_ack <= #1 0;
									multiplier_19_state <= #1 multiplier_19_get_z;
									multiplier_19_input_a_stb <= #1 0;
								end
							end
							multiplier_19_get_z : begin
								if (multiplier_19_output_z_stb) begin
									_r7 <= #1 multiplier_19_output_z;
									multiplier_19_output_z_ack <= #1 1;
									multiplier_19_state <= #1 multiplier_19_put_a;
									multiplier_19_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_19 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_19 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p1rom(input [4:0] rom_bus, output [7:0] rom_value);
	reg [7:0] _rom [0:31];
	initial
	begin
	_rom[0] = 8'b00100000;
	_rom[1] = 8'b00101000;
	_rom[2] = 8'b01010000;
	_rom[3] = 8'b01011001;
	_rom[4] = 8'b00000100;
	_rom[5] = 8'b00001110;
	_rom[6] = 8'b01010010;
	_rom[7] = 8'b01011011;
	_rom[8] = 8'b00000100;
	_rom[9] = 8'b00001110;
	_rom[10] = 8'b01010100;
	_rom[11] = 8'b01011101;
	_rom[12] = 8'b00000100;
	_rom[13] = 8'b00001110;
	_rom[14] = 8'b01010110;
	_rom[15] = 8'b01011111;
	_rom[16] = 8'b00000100;
	_rom[17] = 8'b00001110;
	_rom[18] = 8'b10000000;
	_rom[19] = 8'b10001100;
	_rom[20] = 8'b01100000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p1(clock_signal, reset_signal, rom_bus, rom_value, i0, i0_valid, i0_received, i1, i1_valid, i1_received, i2, i2_valid, i2_received, i3, i3_valid, i3_received, i4, i4_valid, i4_received, i5, i5_valid, i5_received, i6, i6_valid, i6_received, i7, i7_valid, i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [7:0] rom_value;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=3'b000,          // Register addf
			CLR=3'b001,          // Clear register
			I2RW=3'b010,          // Input to register
			J=3'b011,          // Jump to a program location
			R2OWA=3'b100;          // Register to output

	localparam	R0=2'b00,		// Registers in the intructions
			R1=2'b01,
			R2=2'b10,
			R3=2'b11;
	localparam			I0=3'b000,
			I1=3'b001,
			I2=3'b010,
			I3=3'b011,
			I4=3'b100,
			I5=3'b101,
			I6=3'b110,
			I7=3'b111;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:0];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;

	wire [7:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_1_input_a;
	reg [31:0] adder_1_input_b;
	reg adder_1_input_a_stb;
	reg adder_1_input_b_stb;
	reg adder_1_output_z_ack;

	wire [31:0] adder_1_output_z;
	wire adder_1_output_z_stb;
	wire adder_1_input_a_ack;
	wire adder_1_input_b_ack;

	reg	[1:0] adder_1_state;
parameter adder_1_put_a         = 2'd0,
          adder_1_put_b         = 2'd1,
          adder_1_get_z         = 2'd2;
	adder_1 adder_1_inst (adder_1_input_a, adder_1_input_b, adder_1_input_a_stb, adder_1_input_b_stb, adder_1_output_z_ack, clock_signal, reset_signal, adder_1_output_z, adder_1_output_z_stb, adder_1_input_a_ack, adder_1_input_b_ack);


// Start of the component "header" for the opcode clr


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;
	reg i2_recv;
	reg i3_recv;
	reg i4_recv;
	reg i5_recv;
	reg i6_recv;
	reg i7_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i2_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I2 : begin
						if (i2_valid)
						begin
							i2_recv <= #1 1'b1;
						end else begin
							i2_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i2_valid)
						begin
							i2_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i2_valid)
					begin
						i2_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i3_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I3 : begin
						if (i3_valid)
						begin
							i3_recv <= #1 1'b1;
						end else begin
							i3_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i3_valid)
						begin
							i3_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i3_valid)
					begin
						i3_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i4_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I4 : begin
						if (i4_valid)
						begin
							i4_recv <= #1 1'b1;
						end else begin
							i4_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i4_valid)
						begin
							i4_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i4_valid)
					begin
						i4_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i5_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I5 : begin
						if (i5_valid)
						begin
							i5_recv <= #1 1'b1;
						end else begin
							i5_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i5_valid)
						begin
							i5_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i5_valid)
					begin
						i5_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i6_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I6 : begin
						if (i6_valid)
						begin
							i6_recv <= #1 1'b1;
						end else begin
							i6_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i6_valid)
						begin
							i6_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i6_valid)
					begin
						i6_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i7_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I7 : begin
						if (i7_valid)
						begin
							i7_recv <= #1 1'b1;
						end else begin
							i7_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i7_valid)
						begin
							i7_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i7_valid)
					begin
						i7_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				R2OWA: begin
					case (current_instruction[2])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				R2OWA: begin
					case (current_instruction[2])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode clr


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode r2owa

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b ", _r0, _r1, _r2, _r3);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode clr


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode r2owa


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode clr


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode r2owa

				case(current_instruction[7:5])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2:1])
							R2 : begin
							case (adder_1_state)
							adder_1_put_a : begin
								if (adder_1_input_a_ack) begin
									adder_1_input_a <= #1 _r0;
									adder_1_input_a_stb <= #1 1;
									adder_1_output_z_ack <= #1 0;
									adder_1_state <= #1 adder_1_put_b;
								end
							end
							adder_1_put_b : begin
								if (adder_1_input_b_ack) begin
									adder_1_input_b <= #1 _r2;
									adder_1_input_b_stb <= #1 1;
									adder_1_output_z_ack <= #1 0;
									adder_1_state <= #1 adder_1_get_z;
									adder_1_input_a_stb <= #1 0;
								end
							end
							adder_1_get_z : begin
								if (adder_1_output_z_stb) begin
									_r0 <= #1 adder_1_output_z;
									adder_1_output_z_ack <= #1 1;
									adder_1_state <= #1 adder_1_put_a;
									adder_1_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R2");
							end
							R3 : begin
							case (adder_1_state)
							adder_1_put_a : begin
								if (adder_1_input_a_ack) begin
									adder_1_input_a <= #1 _r0;
									adder_1_input_a_stb <= #1 1;
									adder_1_output_z_ack <= #1 0;
									adder_1_state <= #1 adder_1_put_b;
								end
							end
							adder_1_put_b : begin
								if (adder_1_input_b_ack) begin
									adder_1_input_b <= #1 _r3;
									adder_1_input_b_stb <= #1 1;
									adder_1_output_z_ack <= #1 0;
									adder_1_state <= #1 adder_1_get_z;
									adder_1_input_a_stb <= #1 0;
								end
							end
							adder_1_get_z : begin
								if (adder_1_output_z_stb) begin
									_r0 <= #1 adder_1_output_z;
									adder_1_output_z_ack <= #1 1;
									adder_1_state <= #1 adder_1_put_a;
									adder_1_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2:1])
							R2 : begin
							case (adder_1_state)
							adder_1_put_a : begin
								if (adder_1_input_a_ack) begin
									adder_1_input_a <= #1 _r1;
									adder_1_input_a_stb <= #1 1;
									adder_1_output_z_ack <= #1 0;
									adder_1_state <= #1 adder_1_put_b;
								end
							end
							adder_1_put_b : begin
								if (adder_1_input_b_ack) begin
									adder_1_input_b <= #1 _r2;
									adder_1_input_b_stb <= #1 1;
									adder_1_output_z_ack <= #1 0;
									adder_1_state <= #1 adder_1_get_z;
									adder_1_input_a_stb <= #1 0;
								end
							end
							adder_1_get_z : begin
								if (adder_1_output_z_stb) begin
									_r1 <= #1 adder_1_output_z;
									adder_1_output_z_ack <= #1 1;
									adder_1_state <= #1 adder_1_put_a;
									adder_1_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R1 R2");
							end
							R3 : begin
							case (adder_1_state)
							adder_1_put_a : begin
								if (adder_1_input_a_ack) begin
									adder_1_input_a <= #1 _r1;
									adder_1_input_a_stb <= #1 1;
									adder_1_output_z_ack <= #1 0;
									adder_1_state <= #1 adder_1_put_b;
								end
							end
							adder_1_put_b : begin
								if (adder_1_input_b_ack) begin
									adder_1_input_b <= #1 _r3;
									adder_1_input_b_stb <= #1 1;
									adder_1_output_z_ack <= #1 0;
									adder_1_state <= #1 adder_1_get_z;
									adder_1_input_a_stb <= #1 0;
								end
							end
							adder_1_get_z : begin
								if (adder_1_output_z_stb) begin
									_r1 <= #1 adder_1_output_z;
									adder_1_output_z_ack <= #1 1;
									adder_1_state <= #1 adder_1_put_a;
									adder_1_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R1 R3");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode clr

					CLR: begin
						case (current_instruction[4:3])
						R0 : begin
							_r0 <= #1 'b0;
							$display("CLR R0");
						end
						R1 : begin
							_r1 <= #1 'b0;
							$display("CLR R1");
						end
						R2 : begin
							_r2 <= #1 'b0;
							$display("CLR R2");
						end
						R3 : begin
							_r3 <= #1 'b0;
							$display("CLR R3");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r0 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r0 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r0 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r0 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r0 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r0 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I7");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r1 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r1 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r1 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r1 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r1 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r1 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I7");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r2 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r2 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r2 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r2 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r2 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r2 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I7");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r3 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r3 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r3 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r3 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r3 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r3 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I7");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[4:0];
						$display("J ", current_instruction[4:0]);
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						endcase
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign i2_received = i2_recv;
	assign i3_received = i3_recv;
	assign i4_received = i4_recv;
	assign i5_received = i5_recv;
	assign i6_received = i6_recv;
	assign i7_received = i7_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_1 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p20ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b10111111001101010000010011110011;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p20rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p20(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_20_input_a;
	reg [31:0] adder_20_input_b;
	reg adder_20_input_a_stb;
	reg adder_20_input_b_stb;
	reg adder_20_output_z_ack;

	wire [31:0] adder_20_output_z;
	wire adder_20_output_z_stb;
	wire adder_20_input_a_ack;
	wire adder_20_input_b_ack;

	reg	[1:0] adder_20_state;
parameter adder_20_put_a         = 2'd0,
          adder_20_put_b         = 2'd1,
          adder_20_get_z         = 2'd2;
	adder_20 adder_20_inst (adder_20_input_a, adder_20_input_b, adder_20_input_a_stb, adder_20_input_b_stb, adder_20_output_z_ack, clock_signal, reset_signal, adder_20_output_z, adder_20_output_z_stb, adder_20_input_a_ack, adder_20_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_20_input_a;
	reg [31:0] multiplier_20_input_b;
	reg multiplier_20_input_a_stb;
	reg multiplier_20_input_b_stb;
	reg multiplier_20_output_z_ack;

	wire [31:0] multiplier_20_output_z;
	wire multiplier_20_output_z_stb;
	wire multiplier_20_input_a_ack;
	wire multiplier_20_input_b_ack;

	reg	[1:0] multiplier_20_state;
parameter multiplier_20_put_a         = 2'd0,
          multiplier_20_put_b         = 2'd1,
          multiplier_20_get_z         = 2'd2;
	multiplier_20 multiplier_20_inst (multiplier_20_input_a, multiplier_20_input_b, multiplier_20_input_a_stb, multiplier_20_input_b_stb, multiplier_20_output_z_ack, clock_signal, reset_signal, multiplier_20_output_z, multiplier_20_output_z_stb, multiplier_20_input_a_ack, multiplier_20_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_20_state)
							adder_20_put_a : begin
								if (adder_20_input_a_ack) begin
									adder_20_input_a <= #1 _r0;
									adder_20_input_a_stb <= #1 1;
									adder_20_output_z_ack <= #1 0;
									adder_20_state <= #1 adder_20_put_b;
								end
							end
							adder_20_put_b : begin
								if (adder_20_input_b_ack) begin
									adder_20_input_b <= #1 _r7;
									adder_20_input_b_stb <= #1 1;
									adder_20_output_z_ack <= #1 0;
									adder_20_state <= #1 adder_20_get_z;
									adder_20_input_a_stb <= #1 0;
								end
							end
							adder_20_get_z : begin
								if (adder_20_output_z_stb) begin
									_r0 <= #1 adder_20_output_z;
									adder_20_output_z_ack <= #1 1;
									adder_20_state <= #1 adder_20_put_a;
									adder_20_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_20_state)
							adder_20_put_a : begin
								if (adder_20_input_a_ack) begin
									adder_20_input_a <= #1 _r6;
									adder_20_input_a_stb <= #1 1;
									adder_20_output_z_ack <= #1 0;
									adder_20_state <= #1 adder_20_put_b;
								end
							end
							adder_20_put_b : begin
								if (adder_20_input_b_ack) begin
									adder_20_input_b <= #1 _r7;
									adder_20_input_b_stb <= #1 1;
									adder_20_output_z_ack <= #1 0;
									adder_20_state <= #1 adder_20_get_z;
									adder_20_input_a_stb <= #1 0;
								end
							end
							adder_20_get_z : begin
								if (adder_20_output_z_stb) begin
									_r6 <= #1 adder_20_output_z;
									adder_20_output_z_ack <= #1 1;
									adder_20_state <= #1 adder_20_put_a;
									adder_20_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_20_state)
							multiplier_20_put_a : begin
								if (multiplier_20_input_a_ack) begin
									multiplier_20_input_a <= #1 _r0;
									multiplier_20_input_a_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_put_b;
								end
							end
							multiplier_20_put_b : begin
								if (multiplier_20_input_b_ack) begin
									multiplier_20_input_b <= #1 _r3;
									multiplier_20_input_b_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_get_z;
									multiplier_20_input_a_stb <= #1 0;
								end
							end
							multiplier_20_get_z : begin
								if (multiplier_20_output_z_stb) begin
									_r0 <= #1 multiplier_20_output_z;
									multiplier_20_output_z_ack <= #1 1;
									multiplier_20_state <= #1 multiplier_20_put_a;
									multiplier_20_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_20_state)
							multiplier_20_put_a : begin
								if (multiplier_20_input_a_ack) begin
									multiplier_20_input_a <= #1 _r0;
									multiplier_20_input_a_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_put_b;
								end
							end
							multiplier_20_put_b : begin
								if (multiplier_20_input_b_ack) begin
									multiplier_20_input_b <= #1 _r4;
									multiplier_20_input_b_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_get_z;
									multiplier_20_input_a_stb <= #1 0;
								end
							end
							multiplier_20_get_z : begin
								if (multiplier_20_output_z_stb) begin
									_r0 <= #1 multiplier_20_output_z;
									multiplier_20_output_z_ack <= #1 1;
									multiplier_20_state <= #1 multiplier_20_put_a;
									multiplier_20_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_20_state)
							multiplier_20_put_a : begin
								if (multiplier_20_input_a_ack) begin
									multiplier_20_input_a <= #1 _r0;
									multiplier_20_input_a_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_put_b;
								end
							end
							multiplier_20_put_b : begin
								if (multiplier_20_input_b_ack) begin
									multiplier_20_input_b <= #1 _r5;
									multiplier_20_input_b_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_get_z;
									multiplier_20_input_a_stb <= #1 0;
								end
							end
							multiplier_20_get_z : begin
								if (multiplier_20_output_z_stb) begin
									_r0 <= #1 multiplier_20_output_z;
									multiplier_20_output_z_ack <= #1 1;
									multiplier_20_state <= #1 multiplier_20_put_a;
									multiplier_20_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_20_state)
							multiplier_20_put_a : begin
								if (multiplier_20_input_a_ack) begin
									multiplier_20_input_a <= #1 _r7;
									multiplier_20_input_a_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_put_b;
								end
							end
							multiplier_20_put_b : begin
								if (multiplier_20_input_b_ack) begin
									multiplier_20_input_b <= #1 _r3;
									multiplier_20_input_b_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_get_z;
									multiplier_20_input_a_stb <= #1 0;
								end
							end
							multiplier_20_get_z : begin
								if (multiplier_20_output_z_stb) begin
									_r7 <= #1 multiplier_20_output_z;
									multiplier_20_output_z_ack <= #1 1;
									multiplier_20_state <= #1 multiplier_20_put_a;
									multiplier_20_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_20_state)
							multiplier_20_put_a : begin
								if (multiplier_20_input_a_ack) begin
									multiplier_20_input_a <= #1 _r7;
									multiplier_20_input_a_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_put_b;
								end
							end
							multiplier_20_put_b : begin
								if (multiplier_20_input_b_ack) begin
									multiplier_20_input_b <= #1 _r4;
									multiplier_20_input_b_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_get_z;
									multiplier_20_input_a_stb <= #1 0;
								end
							end
							multiplier_20_get_z : begin
								if (multiplier_20_output_z_stb) begin
									_r7 <= #1 multiplier_20_output_z;
									multiplier_20_output_z_ack <= #1 1;
									multiplier_20_state <= #1 multiplier_20_put_a;
									multiplier_20_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_20_state)
							multiplier_20_put_a : begin
								if (multiplier_20_input_a_ack) begin
									multiplier_20_input_a <= #1 _r7;
									multiplier_20_input_a_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_put_b;
								end
							end
							multiplier_20_put_b : begin
								if (multiplier_20_input_b_ack) begin
									multiplier_20_input_b <= #1 _r5;
									multiplier_20_input_b_stb <= #1 1;
									multiplier_20_output_z_ack <= #1 0;
									multiplier_20_state <= #1 multiplier_20_get_z;
									multiplier_20_input_a_stb <= #1 0;
								end
							end
							multiplier_20_get_z : begin
								if (multiplier_20_output_z_stb) begin
									_r7 <= #1 multiplier_20_output_z;
									multiplier_20_output_z_ack <= #1 1;
									multiplier_20_state <= #1 multiplier_20_put_a;
									multiplier_20_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_20 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_20 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p2rom(input [4:0] rom_bus, output [7:0] rom_value);
	reg [7:0] _rom [0:31];
	initial
	begin
	_rom[0] = 8'b00100000;
	_rom[1] = 8'b00101000;
	_rom[2] = 8'b01010000;
	_rom[3] = 8'b01011001;
	_rom[4] = 8'b00000100;
	_rom[5] = 8'b00001110;
	_rom[6] = 8'b01010010;
	_rom[7] = 8'b01011011;
	_rom[8] = 8'b00000100;
	_rom[9] = 8'b00001110;
	_rom[10] = 8'b01010100;
	_rom[11] = 8'b01011101;
	_rom[12] = 8'b00000100;
	_rom[13] = 8'b00001110;
	_rom[14] = 8'b01010110;
	_rom[15] = 8'b01011111;
	_rom[16] = 8'b00000100;
	_rom[17] = 8'b00001110;
	_rom[18] = 8'b10000000;
	_rom[19] = 8'b10001100;
	_rom[20] = 8'b01100000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p2(clock_signal, reset_signal, rom_bus, rom_value, i0, i0_valid, i0_received, i1, i1_valid, i1_received, i2, i2_valid, i2_received, i3, i3_valid, i3_received, i4, i4_valid, i4_received, i5, i5_valid, i5_received, i6, i6_valid, i6_received, i7, i7_valid, i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [7:0] rom_value;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=3'b000,          // Register addf
			CLR=3'b001,          // Clear register
			I2RW=3'b010,          // Input to register
			J=3'b011,          // Jump to a program location
			R2OWA=3'b100;          // Register to output

	localparam	R0=2'b00,		// Registers in the intructions
			R1=2'b01,
			R2=2'b10,
			R3=2'b11;
	localparam			I0=3'b000,
			I1=3'b001,
			I2=3'b010,
			I3=3'b011,
			I4=3'b100,
			I5=3'b101,
			I6=3'b110,
			I7=3'b111;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:0];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;

	wire [7:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_2_input_a;
	reg [31:0] adder_2_input_b;
	reg adder_2_input_a_stb;
	reg adder_2_input_b_stb;
	reg adder_2_output_z_ack;

	wire [31:0] adder_2_output_z;
	wire adder_2_output_z_stb;
	wire adder_2_input_a_ack;
	wire adder_2_input_b_ack;

	reg	[1:0] adder_2_state;
parameter adder_2_put_a         = 2'd0,
          adder_2_put_b         = 2'd1,
          adder_2_get_z         = 2'd2;
	adder_2 adder_2_inst (adder_2_input_a, adder_2_input_b, adder_2_input_a_stb, adder_2_input_b_stb, adder_2_output_z_ack, clock_signal, reset_signal, adder_2_output_z, adder_2_output_z_stb, adder_2_input_a_ack, adder_2_input_b_ack);


// Start of the component "header" for the opcode clr


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;
	reg i2_recv;
	reg i3_recv;
	reg i4_recv;
	reg i5_recv;
	reg i6_recv;
	reg i7_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i2_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I2 : begin
						if (i2_valid)
						begin
							i2_recv <= #1 1'b1;
						end else begin
							i2_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i2_valid)
						begin
							i2_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i2_valid)
					begin
						i2_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i3_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I3 : begin
						if (i3_valid)
						begin
							i3_recv <= #1 1'b1;
						end else begin
							i3_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i3_valid)
						begin
							i3_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i3_valid)
					begin
						i3_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i4_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I4 : begin
						if (i4_valid)
						begin
							i4_recv <= #1 1'b1;
						end else begin
							i4_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i4_valid)
						begin
							i4_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i4_valid)
					begin
						i4_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i5_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I5 : begin
						if (i5_valid)
						begin
							i5_recv <= #1 1'b1;
						end else begin
							i5_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i5_valid)
						begin
							i5_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i5_valid)
					begin
						i5_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i6_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I6 : begin
						if (i6_valid)
						begin
							i6_recv <= #1 1'b1;
						end else begin
							i6_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i6_valid)
						begin
							i6_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i6_valid)
					begin
						i6_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i7_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I7 : begin
						if (i7_valid)
						begin
							i7_recv <= #1 1'b1;
						end else begin
							i7_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i7_valid)
						begin
							i7_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i7_valid)
					begin
						i7_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				R2OWA: begin
					case (current_instruction[2])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				R2OWA: begin
					case (current_instruction[2])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode clr


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode r2owa

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b ", _r0, _r1, _r2, _r3);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode clr


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode r2owa


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode clr


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode r2owa

				case(current_instruction[7:5])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2:1])
							R2 : begin
							case (adder_2_state)
							adder_2_put_a : begin
								if (adder_2_input_a_ack) begin
									adder_2_input_a <= #1 _r0;
									adder_2_input_a_stb <= #1 1;
									adder_2_output_z_ack <= #1 0;
									adder_2_state <= #1 adder_2_put_b;
								end
							end
							adder_2_put_b : begin
								if (adder_2_input_b_ack) begin
									adder_2_input_b <= #1 _r2;
									adder_2_input_b_stb <= #1 1;
									adder_2_output_z_ack <= #1 0;
									adder_2_state <= #1 adder_2_get_z;
									adder_2_input_a_stb <= #1 0;
								end
							end
							adder_2_get_z : begin
								if (adder_2_output_z_stb) begin
									_r0 <= #1 adder_2_output_z;
									adder_2_output_z_ack <= #1 1;
									adder_2_state <= #1 adder_2_put_a;
									adder_2_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R2");
							end
							R3 : begin
							case (adder_2_state)
							adder_2_put_a : begin
								if (adder_2_input_a_ack) begin
									adder_2_input_a <= #1 _r0;
									adder_2_input_a_stb <= #1 1;
									adder_2_output_z_ack <= #1 0;
									adder_2_state <= #1 adder_2_put_b;
								end
							end
							adder_2_put_b : begin
								if (adder_2_input_b_ack) begin
									adder_2_input_b <= #1 _r3;
									adder_2_input_b_stb <= #1 1;
									adder_2_output_z_ack <= #1 0;
									adder_2_state <= #1 adder_2_get_z;
									adder_2_input_a_stb <= #1 0;
								end
							end
							adder_2_get_z : begin
								if (adder_2_output_z_stb) begin
									_r0 <= #1 adder_2_output_z;
									adder_2_output_z_ack <= #1 1;
									adder_2_state <= #1 adder_2_put_a;
									adder_2_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2:1])
							R2 : begin
							case (adder_2_state)
							adder_2_put_a : begin
								if (adder_2_input_a_ack) begin
									adder_2_input_a <= #1 _r1;
									adder_2_input_a_stb <= #1 1;
									adder_2_output_z_ack <= #1 0;
									adder_2_state <= #1 adder_2_put_b;
								end
							end
							adder_2_put_b : begin
								if (adder_2_input_b_ack) begin
									adder_2_input_b <= #1 _r2;
									adder_2_input_b_stb <= #1 1;
									adder_2_output_z_ack <= #1 0;
									adder_2_state <= #1 adder_2_get_z;
									adder_2_input_a_stb <= #1 0;
								end
							end
							adder_2_get_z : begin
								if (adder_2_output_z_stb) begin
									_r1 <= #1 adder_2_output_z;
									adder_2_output_z_ack <= #1 1;
									adder_2_state <= #1 adder_2_put_a;
									adder_2_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R1 R2");
							end
							R3 : begin
							case (adder_2_state)
							adder_2_put_a : begin
								if (adder_2_input_a_ack) begin
									adder_2_input_a <= #1 _r1;
									adder_2_input_a_stb <= #1 1;
									adder_2_output_z_ack <= #1 0;
									adder_2_state <= #1 adder_2_put_b;
								end
							end
							adder_2_put_b : begin
								if (adder_2_input_b_ack) begin
									adder_2_input_b <= #1 _r3;
									adder_2_input_b_stb <= #1 1;
									adder_2_output_z_ack <= #1 0;
									adder_2_state <= #1 adder_2_get_z;
									adder_2_input_a_stb <= #1 0;
								end
							end
							adder_2_get_z : begin
								if (adder_2_output_z_stb) begin
									_r1 <= #1 adder_2_output_z;
									adder_2_output_z_ack <= #1 1;
									adder_2_state <= #1 adder_2_put_a;
									adder_2_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R1 R3");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode clr

					CLR: begin
						case (current_instruction[4:3])
						R0 : begin
							_r0 <= #1 'b0;
							$display("CLR R0");
						end
						R1 : begin
							_r1 <= #1 'b0;
							$display("CLR R1");
						end
						R2 : begin
							_r2 <= #1 'b0;
							$display("CLR R2");
						end
						R3 : begin
							_r3 <= #1 'b0;
							$display("CLR R3");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r0 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r0 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r0 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r0 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r0 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r0 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I7");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r1 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r1 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r1 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r1 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r1 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r1 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I7");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r2 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r2 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r2 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r2 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r2 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r2 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I7");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r3 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r3 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r3 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r3 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r3 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r3 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I7");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[4:0];
						$display("J ", current_instruction[4:0]);
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						endcase
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign i2_received = i2_recv;
	assign i3_received = i3_recv;
	assign i4_received = i4_recv;
	assign i5_received = i5_recv;
	assign i6_received = i6_recv;
	assign i7_received = i7_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_2 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p3rom(input [4:0] rom_bus, output [7:0] rom_value);
	reg [7:0] _rom [0:31];
	initial
	begin
	_rom[0] = 8'b00100000;
	_rom[1] = 8'b00101000;
	_rom[2] = 8'b01010000;
	_rom[3] = 8'b01011001;
	_rom[4] = 8'b00000100;
	_rom[5] = 8'b00001110;
	_rom[6] = 8'b01010010;
	_rom[7] = 8'b01011011;
	_rom[8] = 8'b00000100;
	_rom[9] = 8'b00001110;
	_rom[10] = 8'b01010100;
	_rom[11] = 8'b01011101;
	_rom[12] = 8'b00000100;
	_rom[13] = 8'b00001110;
	_rom[14] = 8'b01010110;
	_rom[15] = 8'b01011111;
	_rom[16] = 8'b00000100;
	_rom[17] = 8'b00001110;
	_rom[18] = 8'b10000000;
	_rom[19] = 8'b10001100;
	_rom[20] = 8'b01100000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p3(clock_signal, reset_signal, rom_bus, rom_value, i0, i0_valid, i0_received, i1, i1_valid, i1_received, i2, i2_valid, i2_received, i3, i3_valid, i3_received, i4, i4_valid, i4_received, i5, i5_valid, i5_received, i6, i6_valid, i6_received, i7, i7_valid, i7_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [7:0] rom_value;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=3'b000,          // Register addf
			CLR=3'b001,          // Clear register
			I2RW=3'b010,          // Input to register
			J=3'b011,          // Jump to a program location
			R2OWA=3'b100;          // Register to output

	localparam	R0=2'b00,		// Registers in the intructions
			R1=2'b01,
			R2=2'b10,
			R3=2'b11;
	localparam			I0=3'b000,
			I1=3'b001,
			I2=3'b010,
			I3=3'b011,
			I4=3'b100,
			I5=3'b101,
			I6=3'b110,
			I7=3'b111;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:0];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;

	wire [7:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_3_input_a;
	reg [31:0] adder_3_input_b;
	reg adder_3_input_a_stb;
	reg adder_3_input_b_stb;
	reg adder_3_output_z_ack;

	wire [31:0] adder_3_output_z;
	wire adder_3_output_z_stb;
	wire adder_3_input_a_ack;
	wire adder_3_input_b_ack;

	reg	[1:0] adder_3_state;
parameter adder_3_put_a         = 2'd0,
          adder_3_put_b         = 2'd1,
          adder_3_get_z         = 2'd2;
	adder_3 adder_3_inst (adder_3_input_a, adder_3_input_b, adder_3_input_a_stb, adder_3_input_b_stb, adder_3_output_z_ack, clock_signal, reset_signal, adder_3_output_z, adder_3_output_z_stb, adder_3_input_a_ack, adder_3_input_b_ack);


// Start of the component "header" for the opcode clr


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;
	reg i2_recv;
	reg i3_recv;
	reg i4_recv;
	reg i5_recv;
	reg i6_recv;
	reg i7_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i2_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I2 : begin
						if (i2_valid)
						begin
							i2_recv <= #1 1'b1;
						end else begin
							i2_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i2_valid)
						begin
							i2_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i2_valid)
					begin
						i2_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i3_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I3 : begin
						if (i3_valid)
						begin
							i3_recv <= #1 1'b1;
						end else begin
							i3_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i3_valid)
						begin
							i3_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i3_valid)
					begin
						i3_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i4_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I4 : begin
						if (i4_valid)
						begin
							i4_recv <= #1 1'b1;
						end else begin
							i4_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i4_valid)
						begin
							i4_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i4_valid)
					begin
						i4_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i5_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I5 : begin
						if (i5_valid)
						begin
							i5_recv <= #1 1'b1;
						end else begin
							i5_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i5_valid)
						begin
							i5_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i5_valid)
					begin
						i5_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i6_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I6 : begin
						if (i6_valid)
						begin
							i6_recv <= #1 1'b1;
						end else begin
							i6_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i6_valid)
						begin
							i6_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i6_valid)
					begin
						i6_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i7_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				I2RW: begin
					case (current_instruction[2:0])
					I7 : begin
						if (i7_valid)
						begin
							i7_recv <= #1 1'b1;
						end else begin
							i7_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i7_valid)
						begin
							i7_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i7_valid)
					begin
						i7_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				R2OWA: begin
					case (current_instruction[2])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[7:5])
				R2OWA: begin
					case (current_instruction[2])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode clr


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode r2owa

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b ", _r0, _r1, _r2, _r3);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode clr


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode r2owa


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode clr


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode r2owa

				case(current_instruction[7:5])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2:1])
							R2 : begin
							case (adder_3_state)
							adder_3_put_a : begin
								if (adder_3_input_a_ack) begin
									adder_3_input_a <= #1 _r0;
									adder_3_input_a_stb <= #1 1;
									adder_3_output_z_ack <= #1 0;
									adder_3_state <= #1 adder_3_put_b;
								end
							end
							adder_3_put_b : begin
								if (adder_3_input_b_ack) begin
									adder_3_input_b <= #1 _r2;
									adder_3_input_b_stb <= #1 1;
									adder_3_output_z_ack <= #1 0;
									adder_3_state <= #1 adder_3_get_z;
									adder_3_input_a_stb <= #1 0;
								end
							end
							adder_3_get_z : begin
								if (adder_3_output_z_stb) begin
									_r0 <= #1 adder_3_output_z;
									adder_3_output_z_ack <= #1 1;
									adder_3_state <= #1 adder_3_put_a;
									adder_3_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R2");
							end
							R3 : begin
							case (adder_3_state)
							adder_3_put_a : begin
								if (adder_3_input_a_ack) begin
									adder_3_input_a <= #1 _r0;
									adder_3_input_a_stb <= #1 1;
									adder_3_output_z_ack <= #1 0;
									adder_3_state <= #1 adder_3_put_b;
								end
							end
							adder_3_put_b : begin
								if (adder_3_input_b_ack) begin
									adder_3_input_b <= #1 _r3;
									adder_3_input_b_stb <= #1 1;
									adder_3_output_z_ack <= #1 0;
									adder_3_state <= #1 adder_3_get_z;
									adder_3_input_a_stb <= #1 0;
								end
							end
							adder_3_get_z : begin
								if (adder_3_output_z_stb) begin
									_r0 <= #1 adder_3_output_z;
									adder_3_output_z_ack <= #1 1;
									adder_3_state <= #1 adder_3_put_a;
									adder_3_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2:1])
							R2 : begin
							case (adder_3_state)
							adder_3_put_a : begin
								if (adder_3_input_a_ack) begin
									adder_3_input_a <= #1 _r1;
									adder_3_input_a_stb <= #1 1;
									adder_3_output_z_ack <= #1 0;
									adder_3_state <= #1 adder_3_put_b;
								end
							end
							adder_3_put_b : begin
								if (adder_3_input_b_ack) begin
									adder_3_input_b <= #1 _r2;
									adder_3_input_b_stb <= #1 1;
									adder_3_output_z_ack <= #1 0;
									adder_3_state <= #1 adder_3_get_z;
									adder_3_input_a_stb <= #1 0;
								end
							end
							adder_3_get_z : begin
								if (adder_3_output_z_stb) begin
									_r1 <= #1 adder_3_output_z;
									adder_3_output_z_ack <= #1 1;
									adder_3_state <= #1 adder_3_put_a;
									adder_3_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R1 R2");
							end
							R3 : begin
							case (adder_3_state)
							adder_3_put_a : begin
								if (adder_3_input_a_ack) begin
									adder_3_input_a <= #1 _r1;
									adder_3_input_a_stb <= #1 1;
									adder_3_output_z_ack <= #1 0;
									adder_3_state <= #1 adder_3_put_b;
								end
							end
							adder_3_put_b : begin
								if (adder_3_input_b_ack) begin
									adder_3_input_b <= #1 _r3;
									adder_3_input_b_stb <= #1 1;
									adder_3_output_z_ack <= #1 0;
									adder_3_state <= #1 adder_3_get_z;
									adder_3_input_a_stb <= #1 0;
								end
							end
							adder_3_get_z : begin
								if (adder_3_output_z_stb) begin
									_r1 <= #1 adder_3_output_z;
									adder_3_output_z_ack <= #1 1;
									adder_3_state <= #1 adder_3_put_a;
									adder_3_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R1 R3");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode clr

					CLR: begin
						case (current_instruction[4:3])
						R0 : begin
							_r0 <= #1 'b0;
							$display("CLR R0");
						end
						R1 : begin
							_r1 <= #1 'b0;
							$display("CLR R1");
						end
						R2 : begin
							_r2 <= #1 'b0;
							$display("CLR R2");
						end
						R3 : begin
							_r3 <= #1 'b0;
							$display("CLR R3");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r0 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r0 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r0 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r0 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r0 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r0 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I7");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r1 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r1 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r1 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r1 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r1 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r1 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I7");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r2 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r2 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r2 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r2 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r2 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r2 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I7");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[2:0])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r3 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r3 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r3 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r3 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r3 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r3 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I7");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[4:0];
						$display("J ", current_instruction[4:0]);
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[4:3])
						R0 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[2])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						endcase
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign i2_received = i2_recv;
	assign i3_received = i3_recv;
	assign i4_received = i4_recv;
	assign i5_received = i5_recv;
	assign i6_received = i6_recv;
	assign i7_received = i7_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_3 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p4ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [2:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:7];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00000000000000000000000000000000;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
		mem[4] = 32'b00000000000000000000000000000000;
		mem[5] = 32'b00000000000000000000000000000000;
		mem[6] = 32'b00000000000000000000000000000000;
		mem[7] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p4rom(input [6:0] rom_bus, output [37:0] rom_value);
	reg [37:0] _rom [0:127];
	initial
	begin
	_rom[0] = 38'b00000100000000000000000000000000000000;
	_rom[1] = 38'b00100000000000000000000000000000000000;
	_rom[2] = 38'b01110001000000000000000000000000000000;
	_rom[3] = 38'b00110100000000000000000000000000000000;
	_rom[4] = 38'b00100000010000000000000000000000000000;
	_rom[5] = 38'b01110001000000000000000000000000000000;
	_rom[6] = 38'b00110100000000000000000000000000000000;
	_rom[7] = 38'b00100000100000000000000000000000000000;
	_rom[8] = 38'b01110001000000000000000000000000000000;
	_rom[9] = 38'b00110100000000000000000000000000000000;
	_rom[10] = 38'b00100000110000000000000000000000000000;
	_rom[11] = 38'b01110001000000000000000000000000000000;
	_rom[12] = 38'b00110100000000000000000000000000000000;
	_rom[13] = 38'b00100001000000000000000000000000000000;
	_rom[14] = 38'b01110001000000000000000000000000000000;
	_rom[15] = 38'b00110100000000000000000000000000000000;
	_rom[16] = 38'b00100001010000000000000000000000000000;
	_rom[17] = 38'b01110001000000000000000000000000000000;
	_rom[18] = 38'b00110100000000000000000000000000000000;
	_rom[19] = 38'b00100001100000000000000000000000000000;
	_rom[20] = 38'b01110001000000000000000000000000000000;
	_rom[21] = 38'b00110100000000000000000000000000000000;
	_rom[22] = 38'b00100001110000000000000000000000000000;
	_rom[23] = 38'b01110001000000000000000000000000000000;
	_rom[24] = 38'b00110100000000000000000000000000000000;
	_rom[25] = 38'b10011000000000000000000000000000000010;
	_rom[26] = 38'b01011010011110000000000000000000000000;
	_rom[27] = 38'b00000100000000000000000000000000000000;
	_rom[28] = 38'b01100001000000000000000000000000000000;
	_rom[29] = 38'b10000010000000000000000000000000000000;
	_rom[30] = 38'b00110100000000000000000000000000000000;
	_rom[31] = 38'b01100001000000000000000000000000000000;
	_rom[32] = 38'b10000010010000000000000000000000000000;
	_rom[33] = 38'b00110100000000000000000000000000000000;
	_rom[34] = 38'b01100001000000000000000000000000000000;
	_rom[35] = 38'b10000010100000000000000000000000000000;
	_rom[36] = 38'b00110100000000000000000000000000000000;
	_rom[37] = 38'b01100001000000000000000000000000000000;
	_rom[38] = 38'b10000010110000000000000000000000000000;
	_rom[39] = 38'b00110100000000000000000000000000000000;
	_rom[40] = 38'b01100001000000000000000000000000000000;
	_rom[41] = 38'b10000011000000000000000000000000000000;
	_rom[42] = 38'b00110100000000000000000000000000000000;
	_rom[43] = 38'b01100001000000000000000000000000000000;
	_rom[44] = 38'b10000011010000000000000000000000000000;
	_rom[45] = 38'b00110100000000000000000000000000000000;
	_rom[46] = 38'b01100001000000000000000000000000000000;
	_rom[47] = 38'b10000011100000000000000000000000000000;
	_rom[48] = 38'b00110100000000000000000000000000000000;
	_rom[49] = 38'b01100001000000000000000000000000000000;
	_rom[50] = 38'b10000011110000000000000000000000000000;
	_rom[51] = 38'b00110100000000000000000000000000000000;
	_rom[52] = 38'b00000100000000000000000000000000000000;
	_rom[53] = 38'b00100010000000000000000000000000000000;
	_rom[54] = 38'b01110001000000000000000000000000000000;
	_rom[55] = 38'b00110100000000000000000000000000000000;
	_rom[56] = 38'b00100010010000000000000000000000000000;
	_rom[57] = 38'b01110001000000000000000000000000000000;
	_rom[58] = 38'b00110100000000000000000000000000000000;
	_rom[59] = 38'b00100010100000000000000000000000000000;
	_rom[60] = 38'b01110001000000000000000000000000000000;
	_rom[61] = 38'b00110100000000000000000000000000000000;
	_rom[62] = 38'b00100010110000000000000000000000000000;
	_rom[63] = 38'b01110001000000000000000000000000000000;
	_rom[64] = 38'b00110100000000000000000000000000000000;
	_rom[65] = 38'b00100011000000000000000000000000000000;
	_rom[66] = 38'b01110001000000000000000000000000000000;
	_rom[67] = 38'b00110100000000000000000000000000000000;
	_rom[68] = 38'b00100011010000000000000000000000000000;
	_rom[69] = 38'b01110001000000000000000000000000000000;
	_rom[70] = 38'b00110100000000000000000000000000000000;
	_rom[71] = 38'b00100011100000000000000000000000000000;
	_rom[72] = 38'b01110001000000000000000000000000000000;
	_rom[73] = 38'b00110100000000000000000000000000000000;
	_rom[74] = 38'b00100011110000000000000000000000000000;
	_rom[75] = 38'b01110001000000000000000000000000000000;
	_rom[76] = 38'b00110100000000000000000000000000000000;
	_rom[77] = 38'b00011000000000000000000000000000000000;
	_rom[78] = 38'b01000011010000000000000000000000000000;
	_rom[79] = 38'b00000100000000000000000000000000000000;
	_rom[80] = 38'b01100001000000000000000000000000000000;
	_rom[81] = 38'b10000000000000000000000000000000000000;
	_rom[82] = 38'b00110100000000000000000000000000000000;
	_rom[83] = 38'b01100001000000000000000000000000000000;
	_rom[84] = 38'b10000000010000000000000000000000000000;
	_rom[85] = 38'b00110100000000000000000000000000000000;
	_rom[86] = 38'b01100001000000000000000000000000000000;
	_rom[87] = 38'b10000000100000000000000000000000000000;
	_rom[88] = 38'b00110100000000000000000000000000000000;
	_rom[89] = 38'b01100001000000000000000000000000000000;
	_rom[90] = 38'b10000000110000000000000000000000000000;
	_rom[91] = 38'b00110100000000000000000000000000000000;
	_rom[92] = 38'b01100001000000000000000000000000000000;
	_rom[93] = 38'b10000001000000000000000000000000000000;
	_rom[94] = 38'b00110100000000000000000000000000000000;
	_rom[95] = 38'b01100001000000000000000000000000000000;
	_rom[96] = 38'b10000001010000000000000000000000000000;
	_rom[97] = 38'b00110100000000000000000000000000000000;
	_rom[98] = 38'b01100001000000000000000000000000000000;
	_rom[99] = 38'b10000001100000000000000000000000000000;
	_rom[100] = 38'b00110100000000000000000000000000000000;
	_rom[101] = 38'b01100001000000000000000000000000000000;
	_rom[102] = 38'b10000001110000000000000000000000000000;
	_rom[103] = 38'b00110100000000000000000000000000000000;
	_rom[104] = 38'b01000000000000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p4(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, i2, i2_valid, i2_received, i3, i3_valid, i3_received, i4, i4_valid, i4_received, i5, i5_valid, i5_received, i6, i6_valid, i6_received, i7, i7_valid, i7_received, i8, i8_valid, i8_received, i9, i9_valid, i9_received, i10, i10_valid, i10_received, i11, i11_valid, i11_received, i12, i12_valid, i12_received, i13, i13_valid, i13_received, i14, i14_valid, i14_received, i15, i15_valid, i15_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received, o2, o2_valid, o2_received, o3, o3_valid, o3_received, o4, o4_valid, o4_received, o5, o5_valid, o5_received, o6, o6_valid, o6_received, o7, o7_valid, o7_received, o8, o8_valid, o8_received, o9, o9_valid, o9_received, o10, o10_valid, o10_received, o11, o11_valid, o11_received, o12, o12_valid, o12_received, o13, o13_valid, o13_received, o14, o14_valid, o14_received, o15, o15_valid, o15_received);

	input clock_signal;
	input reset_signal;
	output  [6:0] rom_bus;
	input  [37:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [2:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	input [31:0] i2;
	input i2_valid;
	output i2_received;
	input [31:0] i3;
	input i3_valid;
	output i3_received;
	input [31:0] i4;
	input i4_valid;
	output i4_received;
	input [31:0] i5;
	input i5_valid;
	output i5_received;
	input [31:0] i6;
	input i6_valid;
	output i6_received;
	input [31:0] i7;
	input i7_valid;
	output i7_received;
	input [31:0] i8;
	input i8_valid;
	output i8_received;
	input [31:0] i9;
	input i9_valid;
	output i9_received;
	input [31:0] i10;
	input i10_valid;
	output i10_received;
	input [31:0] i11;
	input i11_valid;
	output i11_received;
	input [31:0] i12;
	input i12_valid;
	output i12_received;
	input [31:0] i13;
	input i13_valid;
	output i13_received;
	input [31:0] i14;
	input i14_valid;
	output i14_received;
	input [31:0] i15;
	input i15_valid;
	output i15_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;
	output [31:0] o2;
	output o2_valid;
	input o2_received;
	output [31:0] o3;
	output o3_valid;
	input o3_received;
	output [31:0] o4;
	output o4_valid;
	input o4_received;
	output [31:0] o5;
	output o5_valid;
	input o5_received;
	output [31:0] o6;
	output o6_valid;
	input o6_received;
	output [31:0] o7;
	output o7_valid;
	input o7_received;
	output [31:0] o8;
	output o8_valid;
	input o8_received;
	output [31:0] o9;
	output o9_valid;
	input o9_received;
	output [31:0] o10;
	output o10_valid;
	input o10_received;
	output [31:0] o11;
	output o11_valid;
	input o11_received;
	output [31:0] o12;
	output o12_valid;
	input o12_received;
	output [31:0] o13;
	output o13_valid;
	input o13_received;
	output [31:0] o14;
	output o14_valid;
	input o14_received;
	output [31:0] o15;
	output o15_valid;
	input o15_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	CLR=4'b0000,          // Clear register
			DEC=4'b0001,          // Decrement a register by 1
			I2RW=4'b0010,          // Input to register
			INC=4'b0011,          // Increment a register by 1
			J=4'b0100,          // Jump to a program location
			JZ=4'b0101,          // Zero conditional jump
			M2RRI=4'b0110,          // ROM to register
			R2MRI=4'b0111,          // Register indirect copy to RAM
			R2OWA=4'b1000,          // Register to output
			RSET=4'b1001;          // Register set value

	localparam	R0=2'b00,		// Registers in the intructions
			R1=2'b01,
			R2=2'b10,
			R3=2'b11;
	localparam			I0=4'b0000,
			I1=4'b0001,
			I2=4'b0010,
			I3=4'b0011,
			I4=4'b0100,
			I5=4'b0101,
			I6=4'b0110,
			I7=4'b0111,
			I8=4'b1000,
			I9=4'b1001,
			I10=4'b1010,
			I11=4'b1011,
			I12=4'b1100,
			I13=4'b1101,
			I14=4'b1110,
			I15=4'b1111;
	localparam			O0=4'b0000,
			O1=4'b0001,
			O2=4'b0010,
			O3=4'b0011,
			O4=4'b0100,
			O5=4'b0101,
			O6=4'b0110,
			O7=4'b0111,
			O8=4'b1000,
			O9=4'b1001,
			O10=4'b1010,
			O11=4'b1011,
			O12=4'b1100,
			O13=4'b1101,
			O14=4'b1110,
			O15=4'b1111;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;
	reg [31:0] _auxo2;
	reg [31:0] _auxo3;
	reg [31:0] _auxo4;
	reg [31:0] _auxo5;
	reg [31:0] _auxo6;
	reg [31:0] _auxo7;
	reg [31:0] _auxo8;
	reg [31:0] _auxo9;
	reg [31:0] _auxo10;
	reg [31:0] _auxo11;
	reg [31:0] _auxo12;
	reg [31:0] _auxo13;
	reg [31:0] _auxo14;
	reg [31:0] _auxo15;

	reg [31:0] _ram [0:7];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [6:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;

	wire [37:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode clr


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;
	reg i2_recv;
	reg i3_recv;
	reg i4_recv;
	reg i5_recv;
	reg i6_recv;
	reg i7_recv;
	reg i8_recv;
	reg i9_recv;
	reg i10_recv;
	reg i11_recv;
	reg i12_recv;
	reg i13_recv;
	reg i14_recv;
	reg i15_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i2_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I2 : begin
						if (i2_valid)
						begin
							i2_recv <= #1 1'b1;
						end else begin
							i2_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i2_valid)
						begin
							i2_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i2_valid)
					begin
						i2_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i3_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I3 : begin
						if (i3_valid)
						begin
							i3_recv <= #1 1'b1;
						end else begin
							i3_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i3_valid)
						begin
							i3_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i3_valid)
					begin
						i3_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i4_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I4 : begin
						if (i4_valid)
						begin
							i4_recv <= #1 1'b1;
						end else begin
							i4_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i4_valid)
						begin
							i4_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i4_valid)
					begin
						i4_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i5_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I5 : begin
						if (i5_valid)
						begin
							i5_recv <= #1 1'b1;
						end else begin
							i5_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i5_valid)
						begin
							i5_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i5_valid)
					begin
						i5_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i6_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I6 : begin
						if (i6_valid)
						begin
							i6_recv <= #1 1'b1;
						end else begin
							i6_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i6_valid)
						begin
							i6_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i6_valid)
					begin
						i6_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i7_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I7 : begin
						if (i7_valid)
						begin
							i7_recv <= #1 1'b1;
						end else begin
							i7_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i7_valid)
						begin
							i7_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i7_valid)
					begin
						i7_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i8_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I8 : begin
						if (i8_valid)
						begin
							i8_recv <= #1 1'b1;
						end else begin
							i8_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i8_valid)
						begin
							i8_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i8_valid)
					begin
						i8_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i9_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I9 : begin
						if (i9_valid)
						begin
							i9_recv <= #1 1'b1;
						end else begin
							i9_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i9_valid)
						begin
							i9_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i9_valid)
					begin
						i9_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i10_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I10 : begin
						if (i10_valid)
						begin
							i10_recv <= #1 1'b1;
						end else begin
							i10_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i10_valid)
						begin
							i10_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i10_valid)
					begin
						i10_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i11_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I11 : begin
						if (i11_valid)
						begin
							i11_recv <= #1 1'b1;
						end else begin
							i11_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i11_valid)
						begin
							i11_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i11_valid)
					begin
						i11_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i12_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I12 : begin
						if (i12_valid)
						begin
							i12_recv <= #1 1'b1;
						end else begin
							i12_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i12_valid)
						begin
							i12_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i12_valid)
					begin
						i12_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i13_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I13 : begin
						if (i13_valid)
						begin
							i13_recv <= #1 1'b1;
						end else begin
							i13_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i13_valid)
						begin
							i13_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i13_valid)
					begin
						i13_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i14_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I14 : begin
						if (i14_valid)
						begin
							i14_recv <= #1 1'b1;
						end else begin
							i14_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i14_valid)
						begin
							i14_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i14_valid)
					begin
						i14_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i15_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				I2RW: begin
					case (current_instruction[31:28])
					I15 : begin
						if (i15_valid)
						begin
							i15_recv <= #1 1'b1;
						end else begin
							i15_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i15_valid)
						begin
							i15_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i15_valid)
					begin
						i15_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [2:0] addr_ram_m2rri;


// Start of the component "header" for the opcode r2mri

	reg [2:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg o2_val;
	reg o3_val;
	reg o4_val;
	reg o5_val;
	reg o6_val;
	reg o7_val;
	reg o8_val;
	reg o9_val;
	reg o10_val;
	reg o11_val;
	reg o12_val;
	reg o13_val;
	reg o14_val;
	reg o15_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o2_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O2 : begin
						if (waitsm == 1'b1) o2_val <= 1'b1;
					end
					default: begin
						if (o2_received)
						begin
							o2_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o2_received)
					begin
						o2_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o3_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O3 : begin
						if (waitsm == 1'b1) o3_val <= 1'b1;
					end
					default: begin
						if (o3_received)
						begin
							o3_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o3_received)
					begin
						o3_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o4_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O4 : begin
						if (waitsm == 1'b1) o4_val <= 1'b1;
					end
					default: begin
						if (o4_received)
						begin
							o4_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o4_received)
					begin
						o4_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o5_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O5 : begin
						if (waitsm == 1'b1) o5_val <= 1'b1;
					end
					default: begin
						if (o5_received)
						begin
							o5_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o5_received)
					begin
						o5_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o6_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O6 : begin
						if (waitsm == 1'b1) o6_val <= 1'b1;
					end
					default: begin
						if (o6_received)
						begin
							o6_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o6_received)
					begin
						o6_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o7_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O7 : begin
						if (waitsm == 1'b1) o7_val <= 1'b1;
					end
					default: begin
						if (o7_received)
						begin
							o7_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o7_received)
					begin
						o7_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o8_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O8 : begin
						if (waitsm == 1'b1) o8_val <= 1'b1;
					end
					default: begin
						if (o8_received)
						begin
							o8_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o8_received)
					begin
						o8_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o9_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O9 : begin
						if (waitsm == 1'b1) o9_val <= 1'b1;
					end
					default: begin
						if (o9_received)
						begin
							o9_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o9_received)
					begin
						o9_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o10_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O10 : begin
						if (waitsm == 1'b1) o10_val <= 1'b1;
					end
					default: begin
						if (o10_received)
						begin
							o10_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o10_received)
					begin
						o10_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o11_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O11 : begin
						if (waitsm == 1'b1) o11_val <= 1'b1;
					end
					default: begin
						if (o11_received)
						begin
							o11_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o11_received)
					begin
						o11_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o12_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O12 : begin
						if (waitsm == 1'b1) o12_val <= 1'b1;
					end
					default: begin
						if (o12_received)
						begin
							o12_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o12_received)
					begin
						o12_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o13_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O13 : begin
						if (waitsm == 1'b1) o13_val <= 1'b1;
					end
					default: begin
						if (o13_received)
						begin
							o13_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o13_received)
					begin
						o13_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o14_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O14 : begin
						if (waitsm == 1'b1) o14_val <= 1'b1;
					end
					default: begin
						if (o14_received)
						begin
							o14_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o14_received)
					begin
						o14_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o15_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[37:34])
				R2OWA: begin
					case (current_instruction[31:28])
					O15 : begin
						if (waitsm == 1'b1) o15_val <= 1'b1;
					end
					default: begin
						if (o15_received)
						begin
							o15_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o15_received)
					begin
						o15_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 7'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;

// Start of the component "reset" for the opcode clr


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b ", _r0, _r1, _r2, _r3);

// Start of the component "internal state" for the opcode clr


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode clr


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[37:34])

// Start of the component of the "state machine" for the opcode clr

					CLR: begin
						case (current_instruction[33:32])
						R0 : begin
							_r0 <= #1 'b0;
							$display("CLR R0");
						end
						R1 : begin
							_r1 <= #1 'b0;
							$display("CLR R1");
						end
						R2 : begin
							_r2 <= #1 'b0;
							$display("CLR R2");
						end
						R3 : begin
							_r3 <= #1 'b0;
							$display("CLR R3");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[33:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[33:32])
						R0 : begin
							case (current_instruction[31:28])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r0 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r0 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r0 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r0 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r0 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r0 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I7");
								end
							end
							I8 : begin
								if (i8_valid)
								begin
									_r0 <= #1 i8;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I8");
								end
							end
							I9 : begin
								if (i9_valid)
								begin
									_r0 <= #1 i9;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I9");
								end
							end
							I10 : begin
								if (i10_valid)
								begin
									_r0 <= #1 i10;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I10");
								end
							end
							I11 : begin
								if (i11_valid)
								begin
									_r0 <= #1 i11;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I11");
								end
							end
							I12 : begin
								if (i12_valid)
								begin
									_r0 <= #1 i12;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I12");
								end
							end
							I13 : begin
								if (i13_valid)
								begin
									_r0 <= #1 i13;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I13");
								end
							end
							I14 : begin
								if (i14_valid)
								begin
									_r0 <= #1 i14;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I14");
								end
							end
							I15 : begin
								if (i15_valid)
								begin
									_r0 <= #1 i15;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I15");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:28])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r1 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r1 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r1 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r1 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r1 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r1 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I7");
								end
							end
							I8 : begin
								if (i8_valid)
								begin
									_r1 <= #1 i8;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I8");
								end
							end
							I9 : begin
								if (i9_valid)
								begin
									_r1 <= #1 i9;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I9");
								end
							end
							I10 : begin
								if (i10_valid)
								begin
									_r1 <= #1 i10;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I10");
								end
							end
							I11 : begin
								if (i11_valid)
								begin
									_r1 <= #1 i11;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I11");
								end
							end
							I12 : begin
								if (i12_valid)
								begin
									_r1 <= #1 i12;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I12");
								end
							end
							I13 : begin
								if (i13_valid)
								begin
									_r1 <= #1 i13;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I13");
								end
							end
							I14 : begin
								if (i14_valid)
								begin
									_r1 <= #1 i14;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I14");
								end
							end
							I15 : begin
								if (i15_valid)
								begin
									_r1 <= #1 i15;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I15");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:28])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r2 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r2 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r2 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r2 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r2 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r2 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I7");
								end
							end
							I8 : begin
								if (i8_valid)
								begin
									_r2 <= #1 i8;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I8");
								end
							end
							I9 : begin
								if (i9_valid)
								begin
									_r2 <= #1 i9;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I9");
								end
							end
							I10 : begin
								if (i10_valid)
								begin
									_r2 <= #1 i10;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I10");
								end
							end
							I11 : begin
								if (i11_valid)
								begin
									_r2 <= #1 i11;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I11");
								end
							end
							I12 : begin
								if (i12_valid)
								begin
									_r2 <= #1 i12;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I12");
								end
							end
							I13 : begin
								if (i13_valid)
								begin
									_r2 <= #1 i13;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I13");
								end
							end
							I14 : begin
								if (i14_valid)
								begin
									_r2 <= #1 i14;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I14");
								end
							end
							I15 : begin
								if (i15_valid)
								begin
									_r2 <= #1 i15;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I15");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:28])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							I2 : begin
								if (i2_valid)
								begin
									_r3 <= #1 i2;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I2");
								end
							end
							I3 : begin
								if (i3_valid)
								begin
									_r3 <= #1 i3;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I3");
								end
							end
							I4 : begin
								if (i4_valid)
								begin
									_r3 <= #1 i4;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I4");
								end
							end
							I5 : begin
								if (i5_valid)
								begin
									_r3 <= #1 i5;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I5");
								end
							end
							I6 : begin
								if (i6_valid)
								begin
									_r3 <= #1 i6;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I6");
								end
							end
							I7 : begin
								if (i7_valid)
								begin
									_r3 <= #1 i7;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I7");
								end
							end
							I8 : begin
								if (i8_valid)
								begin
									_r3 <= #1 i8;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I8");
								end
							end
							I9 : begin
								if (i9_valid)
								begin
									_r3 <= #1 i9;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I9");
								end
							end
							I10 : begin
								if (i10_valid)
								begin
									_r3 <= #1 i10;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I10");
								end
							end
							I11 : begin
								if (i11_valid)
								begin
									_r3 <= #1 i11;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I11");
								end
							end
							I12 : begin
								if (i12_valid)
								begin
									_r3 <= #1 i12;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I12");
								end
							end
							I13 : begin
								if (i13_valid)
								begin
									_r3 <= #1 i13;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I13");
								end
							end
							I14 : begin
								if (i14_valid)
								begin
									_r3 <= #1 i14;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I14");
								end
							end
							I15 : begin
								if (i15_valid)
								begin
									_r3 <= #1 i15;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I15");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[33:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[33:27];
						$display("J ", current_instruction[33:27]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[33:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:25];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[33:32])
						R0 : begin
							case (current_instruction[31:30])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r0 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R0 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[33:32])
								R0 : begin
									case (current_instruction[31:30])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:30])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:30])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:30])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[33:32])
						R0 : begin
							case (current_instruction[31:28])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							O2 : begin
								if (waitsm == 1'b0) begin
									if (!o2_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo2 <= #1 _r0;
									if (o2_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O2");
							end
							O3 : begin
								if (waitsm == 1'b0) begin
									if (!o3_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo3 <= #1 _r0;
									if (o3_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O3");
							end
							O4 : begin
								if (waitsm == 1'b0) begin
									if (!o4_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo4 <= #1 _r0;
									if (o4_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O4");
							end
							O5 : begin
								if (waitsm == 1'b0) begin
									if (!o5_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo5 <= #1 _r0;
									if (o5_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O5");
							end
							O6 : begin
								if (waitsm == 1'b0) begin
									if (!o6_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo6 <= #1 _r0;
									if (o6_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O6");
							end
							O7 : begin
								if (waitsm == 1'b0) begin
									if (!o7_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo7 <= #1 _r0;
									if (o7_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O7");
							end
							O8 : begin
								if (waitsm == 1'b0) begin
									if (!o8_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo8 <= #1 _r0;
									if (o8_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O8");
							end
							O9 : begin
								if (waitsm == 1'b0) begin
									if (!o9_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo9 <= #1 _r0;
									if (o9_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O9");
							end
							O10 : begin
								if (waitsm == 1'b0) begin
									if (!o10_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo10 <= #1 _r0;
									if (o10_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O10");
							end
							O11 : begin
								if (waitsm == 1'b0) begin
									if (!o11_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo11 <= #1 _r0;
									if (o11_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O11");
							end
							O12 : begin
								if (waitsm == 1'b0) begin
									if (!o12_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo12 <= #1 _r0;
									if (o12_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O12");
							end
							O13 : begin
								if (waitsm == 1'b0) begin
									if (!o13_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo13 <= #1 _r0;
									if (o13_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O13");
							end
							O14 : begin
								if (waitsm == 1'b0) begin
									if (!o14_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo14 <= #1 _r0;
									if (o14_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O14");
							end
							O15 : begin
								if (waitsm == 1'b0) begin
									if (!o15_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo15 <= #1 _r0;
									if (o15_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O15");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:28])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							O2 : begin
								if (waitsm == 1'b0) begin
									if (!o2_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo2 <= #1 _r1;
									if (o2_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O2");
							end
							O3 : begin
								if (waitsm == 1'b0) begin
									if (!o3_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo3 <= #1 _r1;
									if (o3_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O3");
							end
							O4 : begin
								if (waitsm == 1'b0) begin
									if (!o4_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo4 <= #1 _r1;
									if (o4_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O4");
							end
							O5 : begin
								if (waitsm == 1'b0) begin
									if (!o5_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo5 <= #1 _r1;
									if (o5_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O5");
							end
							O6 : begin
								if (waitsm == 1'b0) begin
									if (!o6_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo6 <= #1 _r1;
									if (o6_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O6");
							end
							O7 : begin
								if (waitsm == 1'b0) begin
									if (!o7_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo7 <= #1 _r1;
									if (o7_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O7");
							end
							O8 : begin
								if (waitsm == 1'b0) begin
									if (!o8_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo8 <= #1 _r1;
									if (o8_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O8");
							end
							O9 : begin
								if (waitsm == 1'b0) begin
									if (!o9_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo9 <= #1 _r1;
									if (o9_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O9");
							end
							O10 : begin
								if (waitsm == 1'b0) begin
									if (!o10_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo10 <= #1 _r1;
									if (o10_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O10");
							end
							O11 : begin
								if (waitsm == 1'b0) begin
									if (!o11_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo11 <= #1 _r1;
									if (o11_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O11");
							end
							O12 : begin
								if (waitsm == 1'b0) begin
									if (!o12_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo12 <= #1 _r1;
									if (o12_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O12");
							end
							O13 : begin
								if (waitsm == 1'b0) begin
									if (!o13_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo13 <= #1 _r1;
									if (o13_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O13");
							end
							O14 : begin
								if (waitsm == 1'b0) begin
									if (!o14_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo14 <= #1 _r1;
									if (o14_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O14");
							end
							O15 : begin
								if (waitsm == 1'b0) begin
									if (!o15_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo15 <= #1 _r1;
									if (o15_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O15");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:28])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							O2 : begin
								if (waitsm == 1'b0) begin
									if (!o2_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo2 <= #1 _r2;
									if (o2_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O2");
							end
							O3 : begin
								if (waitsm == 1'b0) begin
									if (!o3_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo3 <= #1 _r2;
									if (o3_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O3");
							end
							O4 : begin
								if (waitsm == 1'b0) begin
									if (!o4_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo4 <= #1 _r2;
									if (o4_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O4");
							end
							O5 : begin
								if (waitsm == 1'b0) begin
									if (!o5_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo5 <= #1 _r2;
									if (o5_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O5");
							end
							O6 : begin
								if (waitsm == 1'b0) begin
									if (!o6_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo6 <= #1 _r2;
									if (o6_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O6");
							end
							O7 : begin
								if (waitsm == 1'b0) begin
									if (!o7_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo7 <= #1 _r2;
									if (o7_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O7");
							end
							O8 : begin
								if (waitsm == 1'b0) begin
									if (!o8_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo8 <= #1 _r2;
									if (o8_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O8");
							end
							O9 : begin
								if (waitsm == 1'b0) begin
									if (!o9_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo9 <= #1 _r2;
									if (o9_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O9");
							end
							O10 : begin
								if (waitsm == 1'b0) begin
									if (!o10_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo10 <= #1 _r2;
									if (o10_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O10");
							end
							O11 : begin
								if (waitsm == 1'b0) begin
									if (!o11_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo11 <= #1 _r2;
									if (o11_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O11");
							end
							O12 : begin
								if (waitsm == 1'b0) begin
									if (!o12_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo12 <= #1 _r2;
									if (o12_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O12");
							end
							O13 : begin
								if (waitsm == 1'b0) begin
									if (!o13_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo13 <= #1 _r2;
									if (o13_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O13");
							end
							O14 : begin
								if (waitsm == 1'b0) begin
									if (!o14_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo14 <= #1 _r2;
									if (o14_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O14");
							end
							O15 : begin
								if (waitsm == 1'b0) begin
									if (!o15_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo15 <= #1 _r2;
									if (o15_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O15");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:28])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							O2 : begin
								if (waitsm == 1'b0) begin
									if (!o2_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo2 <= #1 _r3;
									if (o2_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O2");
							end
							O3 : begin
								if (waitsm == 1'b0) begin
									if (!o3_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo3 <= #1 _r3;
									if (o3_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O3");
							end
							O4 : begin
								if (waitsm == 1'b0) begin
									if (!o4_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo4 <= #1 _r3;
									if (o4_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O4");
							end
							O5 : begin
								if (waitsm == 1'b0) begin
									if (!o5_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo5 <= #1 _r3;
									if (o5_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O5");
							end
							O6 : begin
								if (waitsm == 1'b0) begin
									if (!o6_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo6 <= #1 _r3;
									if (o6_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O6");
							end
							O7 : begin
								if (waitsm == 1'b0) begin
									if (!o7_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo7 <= #1 _r3;
									if (o7_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O7");
							end
							O8 : begin
								if (waitsm == 1'b0) begin
									if (!o8_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo8 <= #1 _r3;
									if (o8_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O8");
							end
							O9 : begin
								if (waitsm == 1'b0) begin
									if (!o9_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo9 <= #1 _r3;
									if (o9_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O9");
							end
							O10 : begin
								if (waitsm == 1'b0) begin
									if (!o10_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo10 <= #1 _r3;
									if (o10_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O10");
							end
							O11 : begin
								if (waitsm == 1'b0) begin
									if (!o11_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo11 <= #1 _r3;
									if (o11_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O11");
							end
							O12 : begin
								if (waitsm == 1'b0) begin
									if (!o12_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo12 <= #1 _r3;
									if (o12_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O12");
							end
							O13 : begin
								if (waitsm == 1'b0) begin
									if (!o13_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo13 <= #1 _r3;
									if (o13_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O13");
							end
							O14 : begin
								if (waitsm == 1'b0) begin
									if (!o14_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo14 <= #1 _r3;
									if (o14_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O14");
							end
							O15 : begin
								if (waitsm == 1'b0) begin
									if (!o15_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo15 <= #1 _r3;
									if (o15_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O15");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[33:32])
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[37:34]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign i2_received = i2_recv;
	assign i3_received = i3_recv;
	assign i4_received = i4_recv;
	assign i5_received = i5_recv;
	assign i6_received = i6_recv;
	assign i7_received = i7_recv;
	assign i8_received = i8_recv;
	assign i9_received = i9_recv;
	assign i10_received = i10_recv;
	assign i11_received = i11_recv;
	assign i12_received = i12_recv;
	assign i13_received = i13_recv;
	assign i14_received = i14_recv;
	assign i15_received = i15_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
	assign o2 = _auxo2;
	assign o2_valid = o2_val;
	assign o3 = _auxo3;
	assign o3_valid = o3_val;
	assign o4 = _auxo4;
	assign o4_valid = o4_val;
	assign o5 = _auxo5;
	assign o5_valid = o5_val;
	assign o6 = _auxo6;
	assign o6_valid = o6_val;
	assign o7 = _auxo7;
	assign o7_valid = o7_val;
	assign o8 = _auxo8;
	assign o8_valid = o8_val;
	assign o9 = _auxo9;
	assign o9_valid = o9_val;
	assign o10 = _auxo10;
	assign o10_valid = o10_val;
	assign o11 = _auxo11;
	assign o11_valid = o11_val;
	assign o12 = _auxo12;
	assign o12_valid = o12_val;
	assign o13 = _auxo13;
	assign o13_valid = o13_val;
	assign o14 = _auxo14;
	assign o14_valid = o14_val;
	assign o15 = _auxo15;
	assign o15_valid = o15_val;
endmodule
`timescale 1ns/1ps
module p5ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00111111001101010000010011110011;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00111111100000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p5rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p5(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_5_input_a;
	reg [31:0] adder_5_input_b;
	reg adder_5_input_a_stb;
	reg adder_5_input_b_stb;
	reg adder_5_output_z_ack;

	wire [31:0] adder_5_output_z;
	wire adder_5_output_z_stb;
	wire adder_5_input_a_ack;
	wire adder_5_input_b_ack;

	reg	[1:0] adder_5_state;
parameter adder_5_put_a         = 2'd0,
          adder_5_put_b         = 2'd1,
          adder_5_get_z         = 2'd2;
	adder_5 adder_5_inst (adder_5_input_a, adder_5_input_b, adder_5_input_a_stb, adder_5_input_b_stb, adder_5_output_z_ack, clock_signal, reset_signal, adder_5_output_z, adder_5_output_z_stb, adder_5_input_a_ack, adder_5_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_5_input_a;
	reg [31:0] multiplier_5_input_b;
	reg multiplier_5_input_a_stb;
	reg multiplier_5_input_b_stb;
	reg multiplier_5_output_z_ack;

	wire [31:0] multiplier_5_output_z;
	wire multiplier_5_output_z_stb;
	wire multiplier_5_input_a_ack;
	wire multiplier_5_input_b_ack;

	reg	[1:0] multiplier_5_state;
parameter multiplier_5_put_a         = 2'd0,
          multiplier_5_put_b         = 2'd1,
          multiplier_5_get_z         = 2'd2;
	multiplier_5 multiplier_5_inst (multiplier_5_input_a, multiplier_5_input_b, multiplier_5_input_a_stb, multiplier_5_input_b_stb, multiplier_5_output_z_ack, clock_signal, reset_signal, multiplier_5_output_z, multiplier_5_output_z_stb, multiplier_5_input_a_ack, multiplier_5_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_5_state)
							adder_5_put_a : begin
								if (adder_5_input_a_ack) begin
									adder_5_input_a <= #1 _r0;
									adder_5_input_a_stb <= #1 1;
									adder_5_output_z_ack <= #1 0;
									adder_5_state <= #1 adder_5_put_b;
								end
							end
							adder_5_put_b : begin
								if (adder_5_input_b_ack) begin
									adder_5_input_b <= #1 _r7;
									adder_5_input_b_stb <= #1 1;
									adder_5_output_z_ack <= #1 0;
									adder_5_state <= #1 adder_5_get_z;
									adder_5_input_a_stb <= #1 0;
								end
							end
							adder_5_get_z : begin
								if (adder_5_output_z_stb) begin
									_r0 <= #1 adder_5_output_z;
									adder_5_output_z_ack <= #1 1;
									adder_5_state <= #1 adder_5_put_a;
									adder_5_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_5_state)
							adder_5_put_a : begin
								if (adder_5_input_a_ack) begin
									adder_5_input_a <= #1 _r6;
									adder_5_input_a_stb <= #1 1;
									adder_5_output_z_ack <= #1 0;
									adder_5_state <= #1 adder_5_put_b;
								end
							end
							adder_5_put_b : begin
								if (adder_5_input_b_ack) begin
									adder_5_input_b <= #1 _r7;
									adder_5_input_b_stb <= #1 1;
									adder_5_output_z_ack <= #1 0;
									adder_5_state <= #1 adder_5_get_z;
									adder_5_input_a_stb <= #1 0;
								end
							end
							adder_5_get_z : begin
								if (adder_5_output_z_stb) begin
									_r6 <= #1 adder_5_output_z;
									adder_5_output_z_ack <= #1 1;
									adder_5_state <= #1 adder_5_put_a;
									adder_5_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_5_state)
							multiplier_5_put_a : begin
								if (multiplier_5_input_a_ack) begin
									multiplier_5_input_a <= #1 _r0;
									multiplier_5_input_a_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_put_b;
								end
							end
							multiplier_5_put_b : begin
								if (multiplier_5_input_b_ack) begin
									multiplier_5_input_b <= #1 _r3;
									multiplier_5_input_b_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_get_z;
									multiplier_5_input_a_stb <= #1 0;
								end
							end
							multiplier_5_get_z : begin
								if (multiplier_5_output_z_stb) begin
									_r0 <= #1 multiplier_5_output_z;
									multiplier_5_output_z_ack <= #1 1;
									multiplier_5_state <= #1 multiplier_5_put_a;
									multiplier_5_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_5_state)
							multiplier_5_put_a : begin
								if (multiplier_5_input_a_ack) begin
									multiplier_5_input_a <= #1 _r0;
									multiplier_5_input_a_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_put_b;
								end
							end
							multiplier_5_put_b : begin
								if (multiplier_5_input_b_ack) begin
									multiplier_5_input_b <= #1 _r4;
									multiplier_5_input_b_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_get_z;
									multiplier_5_input_a_stb <= #1 0;
								end
							end
							multiplier_5_get_z : begin
								if (multiplier_5_output_z_stb) begin
									_r0 <= #1 multiplier_5_output_z;
									multiplier_5_output_z_ack <= #1 1;
									multiplier_5_state <= #1 multiplier_5_put_a;
									multiplier_5_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_5_state)
							multiplier_5_put_a : begin
								if (multiplier_5_input_a_ack) begin
									multiplier_5_input_a <= #1 _r0;
									multiplier_5_input_a_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_put_b;
								end
							end
							multiplier_5_put_b : begin
								if (multiplier_5_input_b_ack) begin
									multiplier_5_input_b <= #1 _r5;
									multiplier_5_input_b_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_get_z;
									multiplier_5_input_a_stb <= #1 0;
								end
							end
							multiplier_5_get_z : begin
								if (multiplier_5_output_z_stb) begin
									_r0 <= #1 multiplier_5_output_z;
									multiplier_5_output_z_ack <= #1 1;
									multiplier_5_state <= #1 multiplier_5_put_a;
									multiplier_5_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_5_state)
							multiplier_5_put_a : begin
								if (multiplier_5_input_a_ack) begin
									multiplier_5_input_a <= #1 _r7;
									multiplier_5_input_a_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_put_b;
								end
							end
							multiplier_5_put_b : begin
								if (multiplier_5_input_b_ack) begin
									multiplier_5_input_b <= #1 _r3;
									multiplier_5_input_b_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_get_z;
									multiplier_5_input_a_stb <= #1 0;
								end
							end
							multiplier_5_get_z : begin
								if (multiplier_5_output_z_stb) begin
									_r7 <= #1 multiplier_5_output_z;
									multiplier_5_output_z_ack <= #1 1;
									multiplier_5_state <= #1 multiplier_5_put_a;
									multiplier_5_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_5_state)
							multiplier_5_put_a : begin
								if (multiplier_5_input_a_ack) begin
									multiplier_5_input_a <= #1 _r7;
									multiplier_5_input_a_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_put_b;
								end
							end
							multiplier_5_put_b : begin
								if (multiplier_5_input_b_ack) begin
									multiplier_5_input_b <= #1 _r4;
									multiplier_5_input_b_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_get_z;
									multiplier_5_input_a_stb <= #1 0;
								end
							end
							multiplier_5_get_z : begin
								if (multiplier_5_output_z_stb) begin
									_r7 <= #1 multiplier_5_output_z;
									multiplier_5_output_z_ack <= #1 1;
									multiplier_5_state <= #1 multiplier_5_put_a;
									multiplier_5_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_5_state)
							multiplier_5_put_a : begin
								if (multiplier_5_input_a_ack) begin
									multiplier_5_input_a <= #1 _r7;
									multiplier_5_input_a_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_put_b;
								end
							end
							multiplier_5_put_b : begin
								if (multiplier_5_input_b_ack) begin
									multiplier_5_input_b <= #1 _r5;
									multiplier_5_input_b_stb <= #1 1;
									multiplier_5_output_z_ack <= #1 0;
									multiplier_5_state <= #1 multiplier_5_get_z;
									multiplier_5_input_a_stb <= #1 0;
								end
							end
							multiplier_5_get_z : begin
								if (multiplier_5_output_z_stb) begin
									_r7 <= #1 multiplier_5_output_z;
									multiplier_5_output_z_ack <= #1 1;
									multiplier_5_state <= #1 multiplier_5_put_a;
									multiplier_5_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_5 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_5 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p6ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00000000000000000000000000000000;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p6rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p6(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_6_input_a;
	reg [31:0] adder_6_input_b;
	reg adder_6_input_a_stb;
	reg adder_6_input_b_stb;
	reg adder_6_output_z_ack;

	wire [31:0] adder_6_output_z;
	wire adder_6_output_z_stb;
	wire adder_6_input_a_ack;
	wire adder_6_input_b_ack;

	reg	[1:0] adder_6_state;
parameter adder_6_put_a         = 2'd0,
          adder_6_put_b         = 2'd1,
          adder_6_get_z         = 2'd2;
	adder_6 adder_6_inst (adder_6_input_a, adder_6_input_b, adder_6_input_a_stb, adder_6_input_b_stb, adder_6_output_z_ack, clock_signal, reset_signal, adder_6_output_z, adder_6_output_z_stb, adder_6_input_a_ack, adder_6_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_6_input_a;
	reg [31:0] multiplier_6_input_b;
	reg multiplier_6_input_a_stb;
	reg multiplier_6_input_b_stb;
	reg multiplier_6_output_z_ack;

	wire [31:0] multiplier_6_output_z;
	wire multiplier_6_output_z_stb;
	wire multiplier_6_input_a_ack;
	wire multiplier_6_input_b_ack;

	reg	[1:0] multiplier_6_state;
parameter multiplier_6_put_a         = 2'd0,
          multiplier_6_put_b         = 2'd1,
          multiplier_6_get_z         = 2'd2;
	multiplier_6 multiplier_6_inst (multiplier_6_input_a, multiplier_6_input_b, multiplier_6_input_a_stb, multiplier_6_input_b_stb, multiplier_6_output_z_ack, clock_signal, reset_signal, multiplier_6_output_z, multiplier_6_output_z_stb, multiplier_6_input_a_ack, multiplier_6_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_6_state)
							adder_6_put_a : begin
								if (adder_6_input_a_ack) begin
									adder_6_input_a <= #1 _r0;
									adder_6_input_a_stb <= #1 1;
									adder_6_output_z_ack <= #1 0;
									adder_6_state <= #1 adder_6_put_b;
								end
							end
							adder_6_put_b : begin
								if (adder_6_input_b_ack) begin
									adder_6_input_b <= #1 _r7;
									adder_6_input_b_stb <= #1 1;
									adder_6_output_z_ack <= #1 0;
									adder_6_state <= #1 adder_6_get_z;
									adder_6_input_a_stb <= #1 0;
								end
							end
							adder_6_get_z : begin
								if (adder_6_output_z_stb) begin
									_r0 <= #1 adder_6_output_z;
									adder_6_output_z_ack <= #1 1;
									adder_6_state <= #1 adder_6_put_a;
									adder_6_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_6_state)
							adder_6_put_a : begin
								if (adder_6_input_a_ack) begin
									adder_6_input_a <= #1 _r6;
									adder_6_input_a_stb <= #1 1;
									adder_6_output_z_ack <= #1 0;
									adder_6_state <= #1 adder_6_put_b;
								end
							end
							adder_6_put_b : begin
								if (adder_6_input_b_ack) begin
									adder_6_input_b <= #1 _r7;
									adder_6_input_b_stb <= #1 1;
									adder_6_output_z_ack <= #1 0;
									adder_6_state <= #1 adder_6_get_z;
									adder_6_input_a_stb <= #1 0;
								end
							end
							adder_6_get_z : begin
								if (adder_6_output_z_stb) begin
									_r6 <= #1 adder_6_output_z;
									adder_6_output_z_ack <= #1 1;
									adder_6_state <= #1 adder_6_put_a;
									adder_6_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_6_state)
							multiplier_6_put_a : begin
								if (multiplier_6_input_a_ack) begin
									multiplier_6_input_a <= #1 _r0;
									multiplier_6_input_a_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_put_b;
								end
							end
							multiplier_6_put_b : begin
								if (multiplier_6_input_b_ack) begin
									multiplier_6_input_b <= #1 _r3;
									multiplier_6_input_b_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_get_z;
									multiplier_6_input_a_stb <= #1 0;
								end
							end
							multiplier_6_get_z : begin
								if (multiplier_6_output_z_stb) begin
									_r0 <= #1 multiplier_6_output_z;
									multiplier_6_output_z_ack <= #1 1;
									multiplier_6_state <= #1 multiplier_6_put_a;
									multiplier_6_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_6_state)
							multiplier_6_put_a : begin
								if (multiplier_6_input_a_ack) begin
									multiplier_6_input_a <= #1 _r0;
									multiplier_6_input_a_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_put_b;
								end
							end
							multiplier_6_put_b : begin
								if (multiplier_6_input_b_ack) begin
									multiplier_6_input_b <= #1 _r4;
									multiplier_6_input_b_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_get_z;
									multiplier_6_input_a_stb <= #1 0;
								end
							end
							multiplier_6_get_z : begin
								if (multiplier_6_output_z_stb) begin
									_r0 <= #1 multiplier_6_output_z;
									multiplier_6_output_z_ack <= #1 1;
									multiplier_6_state <= #1 multiplier_6_put_a;
									multiplier_6_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_6_state)
							multiplier_6_put_a : begin
								if (multiplier_6_input_a_ack) begin
									multiplier_6_input_a <= #1 _r0;
									multiplier_6_input_a_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_put_b;
								end
							end
							multiplier_6_put_b : begin
								if (multiplier_6_input_b_ack) begin
									multiplier_6_input_b <= #1 _r5;
									multiplier_6_input_b_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_get_z;
									multiplier_6_input_a_stb <= #1 0;
								end
							end
							multiplier_6_get_z : begin
								if (multiplier_6_output_z_stb) begin
									_r0 <= #1 multiplier_6_output_z;
									multiplier_6_output_z_ack <= #1 1;
									multiplier_6_state <= #1 multiplier_6_put_a;
									multiplier_6_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_6_state)
							multiplier_6_put_a : begin
								if (multiplier_6_input_a_ack) begin
									multiplier_6_input_a <= #1 _r7;
									multiplier_6_input_a_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_put_b;
								end
							end
							multiplier_6_put_b : begin
								if (multiplier_6_input_b_ack) begin
									multiplier_6_input_b <= #1 _r3;
									multiplier_6_input_b_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_get_z;
									multiplier_6_input_a_stb <= #1 0;
								end
							end
							multiplier_6_get_z : begin
								if (multiplier_6_output_z_stb) begin
									_r7 <= #1 multiplier_6_output_z;
									multiplier_6_output_z_ack <= #1 1;
									multiplier_6_state <= #1 multiplier_6_put_a;
									multiplier_6_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_6_state)
							multiplier_6_put_a : begin
								if (multiplier_6_input_a_ack) begin
									multiplier_6_input_a <= #1 _r7;
									multiplier_6_input_a_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_put_b;
								end
							end
							multiplier_6_put_b : begin
								if (multiplier_6_input_b_ack) begin
									multiplier_6_input_b <= #1 _r4;
									multiplier_6_input_b_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_get_z;
									multiplier_6_input_a_stb <= #1 0;
								end
							end
							multiplier_6_get_z : begin
								if (multiplier_6_output_z_stb) begin
									_r7 <= #1 multiplier_6_output_z;
									multiplier_6_output_z_ack <= #1 1;
									multiplier_6_state <= #1 multiplier_6_put_a;
									multiplier_6_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_6_state)
							multiplier_6_put_a : begin
								if (multiplier_6_input_a_ack) begin
									multiplier_6_input_a <= #1 _r7;
									multiplier_6_input_a_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_put_b;
								end
							end
							multiplier_6_put_b : begin
								if (multiplier_6_input_b_ack) begin
									multiplier_6_input_b <= #1 _r5;
									multiplier_6_input_b_stb <= #1 1;
									multiplier_6_output_z_ack <= #1 0;
									multiplier_6_state <= #1 multiplier_6_get_z;
									multiplier_6_input_a_stb <= #1 0;
								end
							end
							multiplier_6_get_z : begin
								if (multiplier_6_output_z_stb) begin
									_r7 <= #1 multiplier_6_output_z;
									multiplier_6_output_z_ack <= #1 1;
									multiplier_6_state <= #1 multiplier_6_put_a;
									multiplier_6_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_6 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_6 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p7ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00111111001101010000010011110011;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p7rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p7(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_7_input_a;
	reg [31:0] adder_7_input_b;
	reg adder_7_input_a_stb;
	reg adder_7_input_b_stb;
	reg adder_7_output_z_ack;

	wire [31:0] adder_7_output_z;
	wire adder_7_output_z_stb;
	wire adder_7_input_a_ack;
	wire adder_7_input_b_ack;

	reg	[1:0] adder_7_state;
parameter adder_7_put_a         = 2'd0,
          adder_7_put_b         = 2'd1,
          adder_7_get_z         = 2'd2;
	adder_7 adder_7_inst (adder_7_input_a, adder_7_input_b, adder_7_input_a_stb, adder_7_input_b_stb, adder_7_output_z_ack, clock_signal, reset_signal, adder_7_output_z, adder_7_output_z_stb, adder_7_input_a_ack, adder_7_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_7_input_a;
	reg [31:0] multiplier_7_input_b;
	reg multiplier_7_input_a_stb;
	reg multiplier_7_input_b_stb;
	reg multiplier_7_output_z_ack;

	wire [31:0] multiplier_7_output_z;
	wire multiplier_7_output_z_stb;
	wire multiplier_7_input_a_ack;
	wire multiplier_7_input_b_ack;

	reg	[1:0] multiplier_7_state;
parameter multiplier_7_put_a         = 2'd0,
          multiplier_7_put_b         = 2'd1,
          multiplier_7_get_z         = 2'd2;
	multiplier_7 multiplier_7_inst (multiplier_7_input_a, multiplier_7_input_b, multiplier_7_input_a_stb, multiplier_7_input_b_stb, multiplier_7_output_z_ack, clock_signal, reset_signal, multiplier_7_output_z, multiplier_7_output_z_stb, multiplier_7_input_a_ack, multiplier_7_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_7_state)
							adder_7_put_a : begin
								if (adder_7_input_a_ack) begin
									adder_7_input_a <= #1 _r0;
									adder_7_input_a_stb <= #1 1;
									adder_7_output_z_ack <= #1 0;
									adder_7_state <= #1 adder_7_put_b;
								end
							end
							adder_7_put_b : begin
								if (adder_7_input_b_ack) begin
									adder_7_input_b <= #1 _r7;
									adder_7_input_b_stb <= #1 1;
									adder_7_output_z_ack <= #1 0;
									adder_7_state <= #1 adder_7_get_z;
									adder_7_input_a_stb <= #1 0;
								end
							end
							adder_7_get_z : begin
								if (adder_7_output_z_stb) begin
									_r0 <= #1 adder_7_output_z;
									adder_7_output_z_ack <= #1 1;
									adder_7_state <= #1 adder_7_put_a;
									adder_7_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_7_state)
							adder_7_put_a : begin
								if (adder_7_input_a_ack) begin
									adder_7_input_a <= #1 _r6;
									adder_7_input_a_stb <= #1 1;
									adder_7_output_z_ack <= #1 0;
									adder_7_state <= #1 adder_7_put_b;
								end
							end
							adder_7_put_b : begin
								if (adder_7_input_b_ack) begin
									adder_7_input_b <= #1 _r7;
									adder_7_input_b_stb <= #1 1;
									adder_7_output_z_ack <= #1 0;
									adder_7_state <= #1 adder_7_get_z;
									adder_7_input_a_stb <= #1 0;
								end
							end
							adder_7_get_z : begin
								if (adder_7_output_z_stb) begin
									_r6 <= #1 adder_7_output_z;
									adder_7_output_z_ack <= #1 1;
									adder_7_state <= #1 adder_7_put_a;
									adder_7_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_7_state)
							multiplier_7_put_a : begin
								if (multiplier_7_input_a_ack) begin
									multiplier_7_input_a <= #1 _r0;
									multiplier_7_input_a_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_put_b;
								end
							end
							multiplier_7_put_b : begin
								if (multiplier_7_input_b_ack) begin
									multiplier_7_input_b <= #1 _r3;
									multiplier_7_input_b_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_get_z;
									multiplier_7_input_a_stb <= #1 0;
								end
							end
							multiplier_7_get_z : begin
								if (multiplier_7_output_z_stb) begin
									_r0 <= #1 multiplier_7_output_z;
									multiplier_7_output_z_ack <= #1 1;
									multiplier_7_state <= #1 multiplier_7_put_a;
									multiplier_7_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_7_state)
							multiplier_7_put_a : begin
								if (multiplier_7_input_a_ack) begin
									multiplier_7_input_a <= #1 _r0;
									multiplier_7_input_a_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_put_b;
								end
							end
							multiplier_7_put_b : begin
								if (multiplier_7_input_b_ack) begin
									multiplier_7_input_b <= #1 _r4;
									multiplier_7_input_b_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_get_z;
									multiplier_7_input_a_stb <= #1 0;
								end
							end
							multiplier_7_get_z : begin
								if (multiplier_7_output_z_stb) begin
									_r0 <= #1 multiplier_7_output_z;
									multiplier_7_output_z_ack <= #1 1;
									multiplier_7_state <= #1 multiplier_7_put_a;
									multiplier_7_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_7_state)
							multiplier_7_put_a : begin
								if (multiplier_7_input_a_ack) begin
									multiplier_7_input_a <= #1 _r0;
									multiplier_7_input_a_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_put_b;
								end
							end
							multiplier_7_put_b : begin
								if (multiplier_7_input_b_ack) begin
									multiplier_7_input_b <= #1 _r5;
									multiplier_7_input_b_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_get_z;
									multiplier_7_input_a_stb <= #1 0;
								end
							end
							multiplier_7_get_z : begin
								if (multiplier_7_output_z_stb) begin
									_r0 <= #1 multiplier_7_output_z;
									multiplier_7_output_z_ack <= #1 1;
									multiplier_7_state <= #1 multiplier_7_put_a;
									multiplier_7_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_7_state)
							multiplier_7_put_a : begin
								if (multiplier_7_input_a_ack) begin
									multiplier_7_input_a <= #1 _r7;
									multiplier_7_input_a_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_put_b;
								end
							end
							multiplier_7_put_b : begin
								if (multiplier_7_input_b_ack) begin
									multiplier_7_input_b <= #1 _r3;
									multiplier_7_input_b_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_get_z;
									multiplier_7_input_a_stb <= #1 0;
								end
							end
							multiplier_7_get_z : begin
								if (multiplier_7_output_z_stb) begin
									_r7 <= #1 multiplier_7_output_z;
									multiplier_7_output_z_ack <= #1 1;
									multiplier_7_state <= #1 multiplier_7_put_a;
									multiplier_7_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_7_state)
							multiplier_7_put_a : begin
								if (multiplier_7_input_a_ack) begin
									multiplier_7_input_a <= #1 _r7;
									multiplier_7_input_a_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_put_b;
								end
							end
							multiplier_7_put_b : begin
								if (multiplier_7_input_b_ack) begin
									multiplier_7_input_b <= #1 _r4;
									multiplier_7_input_b_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_get_z;
									multiplier_7_input_a_stb <= #1 0;
								end
							end
							multiplier_7_get_z : begin
								if (multiplier_7_output_z_stb) begin
									_r7 <= #1 multiplier_7_output_z;
									multiplier_7_output_z_ack <= #1 1;
									multiplier_7_state <= #1 multiplier_7_put_a;
									multiplier_7_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_7_state)
							multiplier_7_put_a : begin
								if (multiplier_7_input_a_ack) begin
									multiplier_7_input_a <= #1 _r7;
									multiplier_7_input_a_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_put_b;
								end
							end
							multiplier_7_put_b : begin
								if (multiplier_7_input_b_ack) begin
									multiplier_7_input_b <= #1 _r5;
									multiplier_7_input_b_stb <= #1 1;
									multiplier_7_output_z_ack <= #1 0;
									multiplier_7_state <= #1 multiplier_7_get_z;
									multiplier_7_input_a_stb <= #1 0;
								end
							end
							multiplier_7_get_z : begin
								if (multiplier_7_output_z_stb) begin
									_r7 <= #1 multiplier_7_output_z;
									multiplier_7_output_z_ack <= #1 1;
									multiplier_7_state <= #1 multiplier_7_put_a;
									multiplier_7_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_7 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_7 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p8ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00000000000000000000000000000000;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p8rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p8(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_8_input_a;
	reg [31:0] adder_8_input_b;
	reg adder_8_input_a_stb;
	reg adder_8_input_b_stb;
	reg adder_8_output_z_ack;

	wire [31:0] adder_8_output_z;
	wire adder_8_output_z_stb;
	wire adder_8_input_a_ack;
	wire adder_8_input_b_ack;

	reg	[1:0] adder_8_state;
parameter adder_8_put_a         = 2'd0,
          adder_8_put_b         = 2'd1,
          adder_8_get_z         = 2'd2;
	adder_8 adder_8_inst (adder_8_input_a, adder_8_input_b, adder_8_input_a_stb, adder_8_input_b_stb, adder_8_output_z_ack, clock_signal, reset_signal, adder_8_output_z, adder_8_output_z_stb, adder_8_input_a_ack, adder_8_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_8_input_a;
	reg [31:0] multiplier_8_input_b;
	reg multiplier_8_input_a_stb;
	reg multiplier_8_input_b_stb;
	reg multiplier_8_output_z_ack;

	wire [31:0] multiplier_8_output_z;
	wire multiplier_8_output_z_stb;
	wire multiplier_8_input_a_ack;
	wire multiplier_8_input_b_ack;

	reg	[1:0] multiplier_8_state;
parameter multiplier_8_put_a         = 2'd0,
          multiplier_8_put_b         = 2'd1,
          multiplier_8_get_z         = 2'd2;
	multiplier_8 multiplier_8_inst (multiplier_8_input_a, multiplier_8_input_b, multiplier_8_input_a_stb, multiplier_8_input_b_stb, multiplier_8_output_z_ack, clock_signal, reset_signal, multiplier_8_output_z, multiplier_8_output_z_stb, multiplier_8_input_a_ack, multiplier_8_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_8_state)
							adder_8_put_a : begin
								if (adder_8_input_a_ack) begin
									adder_8_input_a <= #1 _r0;
									adder_8_input_a_stb <= #1 1;
									adder_8_output_z_ack <= #1 0;
									adder_8_state <= #1 adder_8_put_b;
								end
							end
							adder_8_put_b : begin
								if (adder_8_input_b_ack) begin
									adder_8_input_b <= #1 _r7;
									adder_8_input_b_stb <= #1 1;
									adder_8_output_z_ack <= #1 0;
									adder_8_state <= #1 adder_8_get_z;
									adder_8_input_a_stb <= #1 0;
								end
							end
							adder_8_get_z : begin
								if (adder_8_output_z_stb) begin
									_r0 <= #1 adder_8_output_z;
									adder_8_output_z_ack <= #1 1;
									adder_8_state <= #1 adder_8_put_a;
									adder_8_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_8_state)
							adder_8_put_a : begin
								if (adder_8_input_a_ack) begin
									adder_8_input_a <= #1 _r6;
									adder_8_input_a_stb <= #1 1;
									adder_8_output_z_ack <= #1 0;
									adder_8_state <= #1 adder_8_put_b;
								end
							end
							adder_8_put_b : begin
								if (adder_8_input_b_ack) begin
									adder_8_input_b <= #1 _r7;
									adder_8_input_b_stb <= #1 1;
									adder_8_output_z_ack <= #1 0;
									adder_8_state <= #1 adder_8_get_z;
									adder_8_input_a_stb <= #1 0;
								end
							end
							adder_8_get_z : begin
								if (adder_8_output_z_stb) begin
									_r6 <= #1 adder_8_output_z;
									adder_8_output_z_ack <= #1 1;
									adder_8_state <= #1 adder_8_put_a;
									adder_8_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_8_state)
							multiplier_8_put_a : begin
								if (multiplier_8_input_a_ack) begin
									multiplier_8_input_a <= #1 _r0;
									multiplier_8_input_a_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_put_b;
								end
							end
							multiplier_8_put_b : begin
								if (multiplier_8_input_b_ack) begin
									multiplier_8_input_b <= #1 _r3;
									multiplier_8_input_b_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_get_z;
									multiplier_8_input_a_stb <= #1 0;
								end
							end
							multiplier_8_get_z : begin
								if (multiplier_8_output_z_stb) begin
									_r0 <= #1 multiplier_8_output_z;
									multiplier_8_output_z_ack <= #1 1;
									multiplier_8_state <= #1 multiplier_8_put_a;
									multiplier_8_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_8_state)
							multiplier_8_put_a : begin
								if (multiplier_8_input_a_ack) begin
									multiplier_8_input_a <= #1 _r0;
									multiplier_8_input_a_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_put_b;
								end
							end
							multiplier_8_put_b : begin
								if (multiplier_8_input_b_ack) begin
									multiplier_8_input_b <= #1 _r4;
									multiplier_8_input_b_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_get_z;
									multiplier_8_input_a_stb <= #1 0;
								end
							end
							multiplier_8_get_z : begin
								if (multiplier_8_output_z_stb) begin
									_r0 <= #1 multiplier_8_output_z;
									multiplier_8_output_z_ack <= #1 1;
									multiplier_8_state <= #1 multiplier_8_put_a;
									multiplier_8_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_8_state)
							multiplier_8_put_a : begin
								if (multiplier_8_input_a_ack) begin
									multiplier_8_input_a <= #1 _r0;
									multiplier_8_input_a_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_put_b;
								end
							end
							multiplier_8_put_b : begin
								if (multiplier_8_input_b_ack) begin
									multiplier_8_input_b <= #1 _r5;
									multiplier_8_input_b_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_get_z;
									multiplier_8_input_a_stb <= #1 0;
								end
							end
							multiplier_8_get_z : begin
								if (multiplier_8_output_z_stb) begin
									_r0 <= #1 multiplier_8_output_z;
									multiplier_8_output_z_ack <= #1 1;
									multiplier_8_state <= #1 multiplier_8_put_a;
									multiplier_8_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_8_state)
							multiplier_8_put_a : begin
								if (multiplier_8_input_a_ack) begin
									multiplier_8_input_a <= #1 _r7;
									multiplier_8_input_a_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_put_b;
								end
							end
							multiplier_8_put_b : begin
								if (multiplier_8_input_b_ack) begin
									multiplier_8_input_b <= #1 _r3;
									multiplier_8_input_b_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_get_z;
									multiplier_8_input_a_stb <= #1 0;
								end
							end
							multiplier_8_get_z : begin
								if (multiplier_8_output_z_stb) begin
									_r7 <= #1 multiplier_8_output_z;
									multiplier_8_output_z_ack <= #1 1;
									multiplier_8_state <= #1 multiplier_8_put_a;
									multiplier_8_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_8_state)
							multiplier_8_put_a : begin
								if (multiplier_8_input_a_ack) begin
									multiplier_8_input_a <= #1 _r7;
									multiplier_8_input_a_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_put_b;
								end
							end
							multiplier_8_put_b : begin
								if (multiplier_8_input_b_ack) begin
									multiplier_8_input_b <= #1 _r4;
									multiplier_8_input_b_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_get_z;
									multiplier_8_input_a_stb <= #1 0;
								end
							end
							multiplier_8_get_z : begin
								if (multiplier_8_output_z_stb) begin
									_r7 <= #1 multiplier_8_output_z;
									multiplier_8_output_z_ack <= #1 1;
									multiplier_8_state <= #1 multiplier_8_put_a;
									multiplier_8_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_8_state)
							multiplier_8_put_a : begin
								if (multiplier_8_input_a_ack) begin
									multiplier_8_input_a <= #1 _r7;
									multiplier_8_input_a_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_put_b;
								end
							end
							multiplier_8_put_b : begin
								if (multiplier_8_input_b_ack) begin
									multiplier_8_input_b <= #1 _r5;
									multiplier_8_input_b_stb <= #1 1;
									multiplier_8_output_z_ack <= #1 0;
									multiplier_8_state <= #1 multiplier_8_get_z;
									multiplier_8_input_a_stb <= #1 0;
								end
							end
							multiplier_8_get_z : begin
								if (multiplier_8_output_z_stb) begin
									_r7 <= #1 multiplier_8_output_z;
									multiplier_8_output_z_ack <= #1 1;
									multiplier_8_state <= #1 multiplier_8_put_a;
									multiplier_8_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_8 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_8 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

`timescale 1ns/1ps
module p9ram(clk, rst, din, dout, addr, wren, en);

	//--------------Input Ports-----------------------
	input clk;
	input rst;
	input [1:0] addr;
	input [31:0] din;
	input wren;
	input en;

	//--------------Inout Ports-----------------------
	output [31:0] dout;

	//--------------Reg-------------------------------
	reg [31:0] mem [0:3];

	reg [31:0] dout_i;

	initial begin
		mem[0] = 32'b00000000000000000000000000000000;
		mem[1] = 32'b00000000000000000000000000000000;
		mem[2] = 32'b00000000000000000000000000000000;
		mem[3] = 32'b00000000000000000000000000000000;
	end
	// Memory Write Block  
	// Write Operation we = 1 
	always @ (posedge clk) 
	begin : MEM_WRITE 
		integer k; 
		if (rst)
		begin 
		end 
		else if (wren)
			mem[addr] <= #1 din;
	end 

	// Memory Read Block
	// Read Operation when we = 0 and oe = 1 
	always @ (posedge clk) 
	begin : MEM_READ 
		if (!wren)
			dout_i <= #1 mem[addr];
	end

	assign dout = dout_i;

endmodule 
`timescale 1ns/1ps
module p9rom(input [4:0] rom_bus, output [38:0] rom_value);
	reg [38:0] _rom [0:31];
	initial
	begin
	_rom[0] = 39'b101101000000000000000000000000000000010;
	_rom[1] = 39'b101100100000000000000000000000000000000;
	_rom[2] = 39'b011001000000000000000000000000000000000;
	_rom[3] = 39'b011101100100000000000000000000000000000;
	_rom[4] = 39'b010000100000000000000000000000000000000;
	_rom[5] = 39'b011110000100000000000000000000000000000;
	_rom[6] = 39'b001100000000000000000000000000000000000;
	_rom[7] = 39'b001110110000000000000000000000000000000;
	_rom[8] = 39'b100000001100000000000000000000000000000;
	_rom[9] = 39'b000111000000000000000000000000000000000;
	_rom[10] = 39'b101111110111111100000000000000000000000;
	_rom[11] = 39'b100011110100000000000000000000000000000;
	_rom[12] = 39'b100011110000000000000000000000000000000;
	_rom[13] = 39'b000011011100000000000000000000000000000;
	_rom[14] = 39'b100000010000000000000000000000000000000;
	_rom[15] = 39'b000111101100000000000000000000000000000;
	_rom[16] = 39'b100011110100000000000000000000000000000;
	_rom[17] = 39'b000000011100000000000000000000000000000;
	_rom[18] = 39'b101011000000000000000000000000000000000;
	_rom[19] = 39'b101000010000000000000000000000000000000;
	_rom[20] = 39'b001001000000000000000000000000000000000;
	_rom[21] = 39'b010000100000000000000000000000000000000;
	_rom[22] = 39'b010100010000000000000000000000000000000;
	_rom[23] = 39'b100100000100000000000000000000000000000;
	end
	assign rom_value = _rom[rom_bus];
endmodule
`timescale 1ns/1ps
module p9(clock_signal, reset_signal, rom_bus, rom_value, ram_din, ram_dout, ram_addr, ram_wren, ram_en, i0, i0_valid, i0_received, i1, i1_valid, i1_received, o0, o0_valid, o0_received, o1, o1_valid, o1_received);

	input clock_signal;
	input reset_signal;
	output  [4:0] rom_bus;
	input  [38:0] rom_value;
	input  [31:0] ram_dout;
	output [31:0] ram_din;
	output  [1:0] ram_addr;
	output ram_wren, ram_en;

	input [31:0] i0;
	input i0_valid;
	output i0_received;
	input [31:0] i1;
	input i1_valid;
	output i1_received;
	output [31:0] o0;
	output o0_valid;
	input o0_received;
	output [31:0] o1;
	output o1_valid;
	input o1_received;

			// Opcodes in the instructions, length according the number of the selected.
	localparam	ADDF=4'b0000,          // Register addf
			CPY=4'b0001,          // Copy from a register to another
			DEC=4'b0010,          // Decrement a register by 1
			I2RW=4'b0011,          // Input to register
			INC=4'b0100,          // Increment a register by 1
			J=4'b0101,          // Jump to a program location
			JZ=4'b0110,          // Zero conditional jump
			M2RRI=4'b0111,          // ROM to register
			MULTF=4'b1000,          // Register float32 multiplcation
			R2MRI=4'b1001,          // Register indirect copy to RAM
			R2OWA=4'b1010,          // Register to output
			RSET=4'b1011;          // Register set value

	localparam	R0=3'b000,		// Registers in the intructions
			R1=3'b001,
			R2=3'b010,
			R3=3'b011,
			R4=3'b100,
			R5=3'b101,
			R6=3'b110,
			R7=3'b111;
	localparam			I0=1'b0,
			I1=1'b1;
	localparam			O0=1'b0,
			O1=1'b1;
	reg [31:0] _auxo0;
	reg [31:0] _auxo1;

	reg [31:0] _ram [0:3];		// Internal processor RAM

	(* KEEP = "TRUE" *) reg [4:0] _pc;		// Program counter

	// The number of registers are 2^R, two letters and an underscore as identifier , maximum R=8 and 265 rigisters
	(* KEEP = "TRUE" *) reg [31:0] _r0;
	(* KEEP = "TRUE" *) reg [31:0] _r1;
	(* KEEP = "TRUE" *) reg [31:0] _r2;
	(* KEEP = "TRUE" *) reg [31:0] _r3;
	(* KEEP = "TRUE" *) reg [31:0] _r4;
	(* KEEP = "TRUE" *) reg [31:0] _r5;
	(* KEEP = "TRUE" *) reg [31:0] _r6;
	(* KEEP = "TRUE" *) reg [31:0] _r7;

	wire [38:0] current_instruction;
	assign current_instruction=rom_value;


// Start of the component "header" for the opcode addf

	reg [31:0] adder_9_input_a;
	reg [31:0] adder_9_input_b;
	reg adder_9_input_a_stb;
	reg adder_9_input_b_stb;
	reg adder_9_output_z_ack;

	wire [31:0] adder_9_output_z;
	wire adder_9_output_z_stb;
	wire adder_9_input_a_ack;
	wire adder_9_input_b_ack;

	reg	[1:0] adder_9_state;
parameter adder_9_put_a         = 2'd0,
          adder_9_put_b         = 2'd1,
          adder_9_get_z         = 2'd2;
	adder_9 adder_9_inst (adder_9_input_a, adder_9_input_b, adder_9_input_a_stb, adder_9_input_b_stb, adder_9_output_z_ack, clock_signal, reset_signal, adder_9_output_z, adder_9_output_z_stb, adder_9_input_a_ack, adder_9_input_b_ack);


// Start of the component "header" for the opcode cpy


// Start of the component "header" for the opcode dec


// Start of the component "header" for the opcode i2rw


	reg i0_recv;
	reg i1_recv;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i0_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I0 : begin
						if (i0_valid)
						begin
							i0_recv <= #1 1'b1;
						end else begin
							i0_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i0_valid)
						begin
							i0_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i0_valid)
					begin
						i0_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			i1_recv <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				I2RW: begin
					case (current_instruction[31])
					I1 : begin
						if (i1_valid)
						begin
							i1_recv <= #1 1'b1;
						end else begin
							i1_recv <= #1 1'b0;
						end
					end
					default: begin
						if (!i1_valid)
						begin
							i1_recv <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (!i1_valid)
					begin
						i1_recv <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode inc


// Start of the component "header" for the opcode j


// Start of the component "header" for the opcode jz


// Start of the component "header" for the opcode m2rri

	//Internal Reg Wire for M2R opcode
	reg state_read_mem_m2rri;
	reg wait_read_mem;
	reg [1:0] addr_ram_m2rri;


// Start of the component "header" for the opcode multf

	reg [31:0] multiplier_9_input_a;
	reg [31:0] multiplier_9_input_b;
	reg multiplier_9_input_a_stb;
	reg multiplier_9_input_b_stb;
	reg multiplier_9_output_z_ack;

	wire [31:0] multiplier_9_output_z;
	wire multiplier_9_output_z_stb;
	wire multiplier_9_input_a_ack;
	wire multiplier_9_input_b_ack;

	reg	[1:0] multiplier_9_state;
parameter multiplier_9_put_a         = 2'd0,
          multiplier_9_put_b         = 2'd1,
          multiplier_9_get_z         = 2'd2;
	multiplier_9 multiplier_9_inst (multiplier_9_input_a, multiplier_9_input_b, multiplier_9_input_a_stb, multiplier_9_input_b_stb, multiplier_9_output_z_ack, clock_signal, reset_signal, multiplier_9_output_z, multiplier_9_output_z_stb, multiplier_9_input_a_ack, multiplier_9_input_b_ack);


// Start of the component "header" for the opcode r2mri

	reg [1:0] addr_ram_to_mem;
	reg [31:0] ram_din_i;
	reg wr_int_ram;

// Start of the component "header" for the opcode r2owa


	reg o0_val;
	reg o1_val;
	reg waitsm;
	initial waitsm = 1'b0;

	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o0_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O0 : begin
						if (waitsm == 1'b1) o0_val <= 1'b1;
					end
					default: begin
						if (o0_received)
						begin
							o0_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o0_received)
					begin
						o0_val <= #1 1'b0;
					end
				end
			endcase
		end
	end
	always @(posedge clock_signal, posedge reset_signal)
	begin
		if (reset_signal)
		begin
			o1_val <= #1 1'b0;
		end
		else
		begin
			case(current_instruction[38:35])
				R2OWA: begin
					case (current_instruction[31])
					O1 : begin
						if (waitsm == 1'b1) o1_val <= 1'b1;
					end
					default: begin
						if (o1_received)
						begin
							o1_val <= #1 1'b0;
						end
					end
					endcase
				end
				default: begin
					if (o1_received)
					begin
						o1_val <= #1 1'b0;
					end
				end
			endcase
		end
	end

// Start of the component "header" for the opcode rset


	always @(posedge clock_signal, posedge reset_signal)
	begin
		if(reset_signal)
		begin
			_pc <= #1 5'h0;
			_r0 <= #1 32'h0;
			_r1 <= #1 32'h0;
			_r2 <= #1 32'h0;
			_r3 <= #1 32'h0;
			_r4 <= #1 32'h0;
			_r5 <= #1 32'h0;
			_r6 <= #1 32'h0;
			_r7 <= #1 32'h0;

// Start of the component "reset" for the opcode addf


// Start of the component "reset" for the opcode cpy


// Start of the component "reset" for the opcode dec


// Start of the component "reset" for the opcode i2rw


// Start of the component "reset" for the opcode inc


// Start of the component "reset" for the opcode j


// Start of the component "reset" for the opcode jz


// Start of the component "reset" for the opcode m2rri


// Start of the component "reset" for the opcode multf


// Start of the component "reset" for the opcode r2mri


// Start of the component "reset" for the opcode r2owa


// Start of the component "reset" for the opcode rset

		end
		else begin
			// ha placeholder
			$display("Program Counter:%d", _pc);
			$display("Instruction:%b", rom_value);
			$display("Registers r0:%b r1:%b r2:%b r3:%b r4:%b r5:%b r6:%b r7:%b ", _r0, _r1, _r2, _r3, _r4, _r5, _r6, _r7);

// Start of the component "internal state" for the opcode addf


// Start of the component "internal state" for the opcode cpy


// Start of the component "internal state" for the opcode dec


// Start of the component "internal state" for the opcode i2rw


// Start of the component "internal state" for the opcode inc


// Start of the component "internal state" for the opcode j


// Start of the component "internal state" for the opcode jz


// Start of the component "internal state" for the opcode m2rri


// Start of the component "internal state" for the opcode multf


// Start of the component "internal state" for the opcode r2mri


// Start of the component "internal state" for the opcode r2owa


// Start of the component "internal state" for the opcode rset


// Start of the component "default state" for the opcode addf


// Start of the component "default state" for the opcode cpy


// Start of the component "default state" for the opcode dec


// Start of the component "default state" for the opcode i2rw


// Start of the component "default state" for the opcode inc


// Start of the component "default state" for the opcode j


// Start of the component "default state" for the opcode jz


// Start of the component "default state" for the opcode m2rri


// Start of the component "default state" for the opcode multf


// Start of the component "default state" for the opcode r2mri


// Start of the component "default state" for the opcode r2owa


// Start of the component "default state" for the opcode rset

				case(current_instruction[38:35])

// Start of the component of the "state machine" for the opcode addf

					ADDF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_9_state)
							adder_9_put_a : begin
								if (adder_9_input_a_ack) begin
									adder_9_input_a <= #1 _r0;
									adder_9_input_a_stb <= #1 1;
									adder_9_output_z_ack <= #1 0;
									adder_9_state <= #1 adder_9_put_b;
								end
							end
							adder_9_put_b : begin
								if (adder_9_input_b_ack) begin
									adder_9_input_b <= #1 _r7;
									adder_9_input_b_stb <= #1 1;
									adder_9_output_z_ack <= #1 0;
									adder_9_state <= #1 adder_9_get_z;
									adder_9_input_a_stb <= #1 0;
								end
							end
							adder_9_get_z : begin
								if (adder_9_output_z_stb) begin
									_r0 <= #1 adder_9_output_z;
									adder_9_output_z_ack <= #1 1;
									adder_9_state <= #1 adder_9_put_a;
									adder_9_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R7 : begin
							case (adder_9_state)
							adder_9_put_a : begin
								if (adder_9_input_a_ack) begin
									adder_9_input_a <= #1 _r6;
									adder_9_input_a_stb <= #1 1;
									adder_9_output_z_ack <= #1 0;
									adder_9_state <= #1 adder_9_put_b;
								end
							end
							adder_9_put_b : begin
								if (adder_9_input_b_ack) begin
									adder_9_input_b <= #1 _r7;
									adder_9_input_b_stb <= #1 1;
									adder_9_output_z_ack <= #1 0;
									adder_9_state <= #1 adder_9_get_z;
									adder_9_input_a_stb <= #1 0;
								end
							end
							adder_9_get_z : begin
								if (adder_9_output_z_stb) begin
									_r6 <= #1 adder_9_output_z;
									adder_9_output_z_ack <= #1 1;
									adder_9_state <= #1 adder_9_put_a;
									adder_9_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R6 R7");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode cpy

					CPY: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r0 <= #1 _r0;
								$display("CPY R0 R0");
							end
							R1 : begin
								_r0 <= #1 _r1;
								$display("CPY R0 R1");
							end
							R2 : begin
								_r0 <= #1 _r2;
								$display("CPY R0 R2");
							end
							R3 : begin
								_r0 <= #1 _r3;
								$display("CPY R0 R3");
							end
							R4 : begin
								_r0 <= #1 _r4;
								$display("CPY R0 R4");
							end
							R5 : begin
								_r0 <= #1 _r5;
								$display("CPY R0 R5");
							end
							R6 : begin
								_r0 <= #1 _r6;
								$display("CPY R0 R6");
							end
							R7 : begin
								_r0 <= #1 _r7;
								$display("CPY R0 R7");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r1 <= #1 _r0;
								$display("CPY R1 R0");
							end
							R1 : begin
								_r1 <= #1 _r1;
								$display("CPY R1 R1");
							end
							R2 : begin
								_r1 <= #1 _r2;
								$display("CPY R1 R2");
							end
							R3 : begin
								_r1 <= #1 _r3;
								$display("CPY R1 R3");
							end
							R4 : begin
								_r1 <= #1 _r4;
								$display("CPY R1 R4");
							end
							R5 : begin
								_r1 <= #1 _r5;
								$display("CPY R1 R5");
							end
							R6 : begin
								_r1 <= #1 _r6;
								$display("CPY R1 R6");
							end
							R7 : begin
								_r1 <= #1 _r7;
								$display("CPY R1 R7");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r2 <= #1 _r0;
								$display("CPY R2 R0");
							end
							R1 : begin
								_r2 <= #1 _r1;
								$display("CPY R2 R1");
							end
							R2 : begin
								_r2 <= #1 _r2;
								$display("CPY R2 R2");
							end
							R3 : begin
								_r2 <= #1 _r3;
								$display("CPY R2 R3");
							end
							R4 : begin
								_r2 <= #1 _r4;
								$display("CPY R2 R4");
							end
							R5 : begin
								_r2 <= #1 _r5;
								$display("CPY R2 R5");
							end
							R6 : begin
								_r2 <= #1 _r6;
								$display("CPY R2 R6");
							end
							R7 : begin
								_r2 <= #1 _r7;
								$display("CPY R2 R7");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r3 <= #1 _r0;
								$display("CPY R3 R0");
							end
							R1 : begin
								_r3 <= #1 _r1;
								$display("CPY R3 R1");
							end
							R2 : begin
								_r3 <= #1 _r2;
								$display("CPY R3 R2");
							end
							R3 : begin
								_r3 <= #1 _r3;
								$display("CPY R3 R3");
							end
							R4 : begin
								_r3 <= #1 _r4;
								$display("CPY R3 R4");
							end
							R5 : begin
								_r3 <= #1 _r5;
								$display("CPY R3 R5");
							end
							R6 : begin
								_r3 <= #1 _r6;
								$display("CPY R3 R6");
							end
							R7 : begin
								_r3 <= #1 _r7;
								$display("CPY R3 R7");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r4 <= #1 _r0;
								$display("CPY R4 R0");
							end
							R1 : begin
								_r4 <= #1 _r1;
								$display("CPY R4 R1");
							end
							R2 : begin
								_r4 <= #1 _r2;
								$display("CPY R4 R2");
							end
							R3 : begin
								_r4 <= #1 _r3;
								$display("CPY R4 R3");
							end
							R4 : begin
								_r4 <= #1 _r4;
								$display("CPY R4 R4");
							end
							R5 : begin
								_r4 <= #1 _r5;
								$display("CPY R4 R5");
							end
							R6 : begin
								_r4 <= #1 _r6;
								$display("CPY R4 R6");
							end
							R7 : begin
								_r4 <= #1 _r7;
								$display("CPY R4 R7");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r5 <= #1 _r0;
								$display("CPY R5 R0");
							end
							R1 : begin
								_r5 <= #1 _r1;
								$display("CPY R5 R1");
							end
							R2 : begin
								_r5 <= #1 _r2;
								$display("CPY R5 R2");
							end
							R3 : begin
								_r5 <= #1 _r3;
								$display("CPY R5 R3");
							end
							R4 : begin
								_r5 <= #1 _r4;
								$display("CPY R5 R4");
							end
							R5 : begin
								_r5 <= #1 _r5;
								$display("CPY R5 R5");
							end
							R6 : begin
								_r5 <= #1 _r6;
								$display("CPY R5 R6");
							end
							R7 : begin
								_r5 <= #1 _r7;
								$display("CPY R5 R7");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r6 <= #1 _r0;
								$display("CPY R6 R0");
							end
							R1 : begin
								_r6 <= #1 _r1;
								$display("CPY R6 R1");
							end
							R2 : begin
								_r6 <= #1 _r2;
								$display("CPY R6 R2");
							end
							R3 : begin
								_r6 <= #1 _r3;
								$display("CPY R6 R3");
							end
							R4 : begin
								_r6 <= #1 _r4;
								$display("CPY R6 R4");
							end
							R5 : begin
								_r6 <= #1 _r5;
								$display("CPY R6 R5");
							end
							R6 : begin
								_r6 <= #1 _r6;
								$display("CPY R6 R6");
							end
							R7 : begin
								_r6 <= #1 _r7;
								$display("CPY R6 R7");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R0 : begin
								_r7 <= #1 _r0;
								$display("CPY R7 R0");
							end
							R1 : begin
								_r7 <= #1 _r1;
								$display("CPY R7 R1");
							end
							R2 : begin
								_r7 <= #1 _r2;
								$display("CPY R7 R2");
							end
							R3 : begin
								_r7 <= #1 _r3;
								$display("CPY R7 R3");
							end
							R4 : begin
								_r7 <= #1 _r4;
								$display("CPY R7 R4");
							end
							R5 : begin
								_r7 <= #1 _r5;
								$display("CPY R7 R5");
							end
							R6 : begin
								_r7 <= #1 _r6;
								$display("CPY R7 R6");
							end
							R7 : begin
								_r7 <= #1 _r7;
								$display("CPY R7 R7");
							end
							endcase
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode dec

					DEC: begin
						case (current_instruction[34:32])
						R2 : begin
							_r2 <= _r2 - 1'b1;
							$display("DEC R2");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode i2rw

					I2RW: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r0 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r0 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R0 I1");
								end
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r1 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r1 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R1 I1");
								end
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r2 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r2 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R2 I1");
								end
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r3 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r3 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R3 I1");
								end
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r4 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r4 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R4 I1");
								end
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r5 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r5 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R5 I1");
								end
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r6 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r6 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R6 I1");
								end
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							I0 : begin
								if (i0_valid)
								begin
									_r7 <= #1 i0;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I0");
								end
							end
							I1 : begin
								if (i1_valid)
								begin
									_r7 <= #1 i1;
									_pc <= #1 _pc + 1'b1;
									$display("I2RW R7 I1");
								end
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode inc

					INC: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 _r1 + 1'b1;
							$display("INC R1");
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end

// Start of the component of the "state machine" for the opcode j

					J: begin
						_pc <= #1 current_instruction[34:30];
						$display("J ", current_instruction[34:30]);
					end

// Start of the component of the "state machine" for the opcode jz

					JZ: begin
						case (current_instruction[34:32])
							R2 : begin
								if(_r2 == 'b0) begin
								_pc <= #1 current_instruction[31:27];
								end
								else begin
									_pc <= #1 _pc + 1'b1;
								end
								$display("JZ R2 ",_r2);
							end
						endcase
					end

// Start of the component of the "state machine" for the opcode m2rri

					M2RRI: begin
						case (current_instruction[34:32])
						R3 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r3 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R3 ",_r1);
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31:29])
							R1 : begin
								if (state_read_mem_m2rri == 1'b1) begin
									_r4 <= #1 ram_dout;
									state_read_mem_m2rri <= 1'b0;
									_pc <= #1 _pc + 1'b1;
								end
								else begin
									if (wait_read_mem == 1'b1) begin
										state_read_mem_m2rri <= 1'b1;
										wait_read_mem <= 1'b0;
									end
									else begin
										wait_read_mem <= 1'b1;
										addr_ram_m2rri <= #1 _r1;
									end
								end
								$display("M2RRI R4 ",_r1);
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode multf

					MULTF: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_9_state)
							multiplier_9_put_a : begin
								if (multiplier_9_input_a_ack) begin
									multiplier_9_input_a <= #1 _r0;
									multiplier_9_input_a_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_put_b;
								end
							end
							multiplier_9_put_b : begin
								if (multiplier_9_input_b_ack) begin
									multiplier_9_input_b <= #1 _r3;
									multiplier_9_input_b_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_get_z;
									multiplier_9_input_a_stb <= #1 0;
								end
							end
							multiplier_9_get_z : begin
								if (multiplier_9_output_z_stb) begin
									_r0 <= #1 multiplier_9_output_z;
									multiplier_9_output_z_ack <= #1 1;
									multiplier_9_state <= #1 multiplier_9_put_a;
									multiplier_9_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R3");
							end
							R4 : begin
							case (multiplier_9_state)
							multiplier_9_put_a : begin
								if (multiplier_9_input_a_ack) begin
									multiplier_9_input_a <= #1 _r0;
									multiplier_9_input_a_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_put_b;
								end
							end
							multiplier_9_put_b : begin
								if (multiplier_9_input_b_ack) begin
									multiplier_9_input_b <= #1 _r4;
									multiplier_9_input_b_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_get_z;
									multiplier_9_input_a_stb <= #1 0;
								end
							end
							multiplier_9_get_z : begin
								if (multiplier_9_output_z_stb) begin
									_r0 <= #1 multiplier_9_output_z;
									multiplier_9_output_z_ack <= #1 1;
									multiplier_9_state <= #1 multiplier_9_put_a;
									multiplier_9_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R4");
							end
							R5 : begin
							case (multiplier_9_state)
							multiplier_9_put_a : begin
								if (multiplier_9_input_a_ack) begin
									multiplier_9_input_a <= #1 _r0;
									multiplier_9_input_a_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_put_b;
								end
							end
							multiplier_9_put_b : begin
								if (multiplier_9_input_b_ack) begin
									multiplier_9_input_b <= #1 _r5;
									multiplier_9_input_b_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_get_z;
									multiplier_9_input_a_stb <= #1 0;
								end
							end
							multiplier_9_get_z : begin
								if (multiplier_9_output_z_stb) begin
									_r0 <= #1 multiplier_9_output_z;
									multiplier_9_output_z_ack <= #1 1;
									multiplier_9_state <= #1 multiplier_9_put_a;
									multiplier_9_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R0 R5");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31:29])
							R3 : begin
							case (multiplier_9_state)
							multiplier_9_put_a : begin
								if (multiplier_9_input_a_ack) begin
									multiplier_9_input_a <= #1 _r7;
									multiplier_9_input_a_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_put_b;
								end
							end
							multiplier_9_put_b : begin
								if (multiplier_9_input_b_ack) begin
									multiplier_9_input_b <= #1 _r3;
									multiplier_9_input_b_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_get_z;
									multiplier_9_input_a_stb <= #1 0;
								end
							end
							multiplier_9_get_z : begin
								if (multiplier_9_output_z_stb) begin
									_r7 <= #1 multiplier_9_output_z;
									multiplier_9_output_z_ack <= #1 1;
									multiplier_9_state <= #1 multiplier_9_put_a;
									multiplier_9_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R3");
							end
							R4 : begin
							case (multiplier_9_state)
							multiplier_9_put_a : begin
								if (multiplier_9_input_a_ack) begin
									multiplier_9_input_a <= #1 _r7;
									multiplier_9_input_a_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_put_b;
								end
							end
							multiplier_9_put_b : begin
								if (multiplier_9_input_b_ack) begin
									multiplier_9_input_b <= #1 _r4;
									multiplier_9_input_b_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_get_z;
									multiplier_9_input_a_stb <= #1 0;
								end
							end
							multiplier_9_get_z : begin
								if (multiplier_9_output_z_stb) begin
									_r7 <= #1 multiplier_9_output_z;
									multiplier_9_output_z_ack <= #1 1;
									multiplier_9_state <= #1 multiplier_9_put_a;
									multiplier_9_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R4");
							end
							R5 : begin
							case (multiplier_9_state)
							multiplier_9_put_a : begin
								if (multiplier_9_input_a_ack) begin
									multiplier_9_input_a <= #1 _r7;
									multiplier_9_input_a_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_put_b;
								end
							end
							multiplier_9_put_b : begin
								if (multiplier_9_input_b_ack) begin
									multiplier_9_input_b <= #1 _r5;
									multiplier_9_input_b_stb <= #1 1;
									multiplier_9_output_z_ack <= #1 0;
									multiplier_9_state <= #1 multiplier_9_get_z;
									multiplier_9_input_a_stb <= #1 0;
								end
							end
							multiplier_9_get_z : begin
								if (multiplier_9_output_z_stb) begin
									_r7 <= #1 multiplier_9_output_z;
									multiplier_9_output_z_ack <= #1 1;
									multiplier_9_state <= #1 multiplier_9_put_a;
									multiplier_9_input_b_stb <= #1 0;
									_pc <= #1 _pc + 1'b1;
								end
							end
							endcase
								$display("ADDF R7 R5");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode r2mri

					R2MRI: begin
						if (wr_int_ram == 0) begin
							wr_int_ram <= #1 1'b1;
							case (current_instruction[34:32])
								R0 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r0;
											$display("R2MRI R0 ",_r7);
										end
									endcase
								end
								R1 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r1;
											$display("R2MRI R1 ",_r7);
										end
									endcase
								end
								R2 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r2;
											$display("R2MRI R2 ",_r7);
										end
									endcase
								end
								R3 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r3;
											$display("R2MRI R3 ",_r7);
										end
									endcase
								end
								R4 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r4;
											$display("R2MRI R4 ",_r7);
										end
									endcase
								end
								R5 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r5;
											$display("R2MRI R5 ",_r7);
										end
									endcase
								end
								R6 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r6;
											$display("R2MRI R6 ",_r7);
										end
									endcase
								end
								R7 : begin
									case (current_instruction[31:29])
										R0 : begin
											addr_ram_to_mem <= _r0;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r0);
										end
										R1 : begin
											addr_ram_to_mem <= _r1;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r1);
										end
										R2 : begin
											addr_ram_to_mem <= _r2;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r2);
										end
										R3 : begin
											addr_ram_to_mem <= _r3;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r3);
										end
										R4 : begin
											addr_ram_to_mem <= _r4;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r4);
										end
										R5 : begin
											addr_ram_to_mem <= _r5;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r5);
										end
										R6 : begin
											addr_ram_to_mem <= _r6;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r6);
										end
										R7 : begin
											addr_ram_to_mem <= _r7;
											ram_din_i <= _r7;
											$display("R2MRI R7 ",_r7);
										end
									endcase
								end
							endcase
						end
						else begin
							wr_int_ram <= #1 1'b0;
							_pc <= #1 _pc + 1'b1;
						end
					end

// Start of the component of the "state machine" for the opcode r2owa

					R2OWA: begin
						case (current_instruction[34:32])
						R0 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r0;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r0;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R0 O1");
							end
							endcase
						end
						R1 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r1;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r1;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R1 O1");
							end
							endcase
						end
						R2 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r2;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r2;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R2 O1");
							end
							endcase
						end
						R3 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r3;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r3;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R3 O1");
							end
							endcase
						end
						R4 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r4;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r4;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R4 O1");
							end
							endcase
						end
						R5 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r5;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r5;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R5 O1");
							end
							endcase
						end
						R6 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r6;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r6;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R6 O1");
							end
							endcase
						end
						R7 : begin
							case (current_instruction[31])
							O0 : begin
								if (waitsm == 1'b0) begin
									if (!o0_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo0 <= #1 _r7;
									if (o0_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O0");
							end
							O1 : begin
								if (waitsm == 1'b0) begin
									if (!o1_received) begin
										waitsm <= 1'b1;
									end
								end else begin
									_auxo1 <= #1 _r7;
									if (o1_received) begin
										_pc <= #1 _pc + 1'b1;
										waitsm <= 1'b0;
									end
								end
								$display("R2OWA R7 O1");
							end
							endcase
						end
						endcase
					end

// Start of the component of the "state machine" for the opcode rset

					RSET: begin
						case (current_instruction[34:32])
						R1 : begin
							_r1 <= #1 current_instruction[31:0];
							$display("RSET R1 ",_r1);
						end
						R2 : begin
							_r2 <= #1 current_instruction[31:0];
							$display("RSET R2 ",_r2);
						end
						R7 : begin
							_r7 <= #1 current_instruction[31:0];
							$display("RSET R7 ",_r7);
						end
						endcase
						_pc <= #1 _pc + 1'b1;
					end
					default : begin
						$display("Unknown Opcode");
						_pc <= #1 _pc + 1'b1;
					end
				endcase
			// ha placeholder
		end
	end
	assign rom_bus = _pc;
	assign ram_en = 1'b1;
	assign ram_addr =  (current_instruction[38:35]==M2RRI) ? addr_ram_m2rri: addr_ram_to_mem;
	assign ram_din = ram_din_i;
	assign ram_wren = wr_int_ram;
	assign i0_received = i0_recv;
	assign i1_received = i1_recv;
	assign o0 = _auxo0;
	assign o0_valid = o0_val;
	assign o1 = _auxo1;
	assign o1_valid = o1_val;
endmodule

//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module adder_9 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            align         = 4'd4,
            add_0         = 4'd5,
            add_1         = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [31:0] a, b, z;
  reg       [26:0] a_m, b_m;
  reg       [23:0] z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [27:0] sum;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= {a[22 : 0], 3'd0};
        b_m <= {b[22 : 0], 3'd0};
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is inf and signs don't match return nan
          if ((b_e == 128) && (a_s != b_s)) begin
              z[31] <= b_s;
              z[30:23] <= 255;
              z[22] <= 1;
              z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          state <= put_z;
        //if a is zero return b
        end else if ((($signed(a_e) == -127) && (a_m == 0)) && (($signed(b_e) == -127) && (b_m == 0))) begin
          z[31] <= a_s & b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if a is zero return b
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= b_s;
          z[30:23] <= b_e[7:0] + 127;
          z[22:0] <= b_m[26:3];
          state <= put_z;
        //if b is zero return a
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s;
          z[30:23] <= a_e[7:0] + 127;
          z[22:0] <= a_m[26:3];
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[26] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[26] <= 1;
          end
          state <= align;
        end
      end

      align:
      begin
        if ($signed(a_e) > $signed(b_e)) begin
          b_e <= b_e + 1;
          b_m <= b_m >> 1;
          b_m[0] <= b_m[0] | b_m[1];
        end else if ($signed(a_e) < $signed(b_e)) begin
          a_e <= a_e + 1;
          a_m <= a_m >> 1;
          a_m[0] <= a_m[0] | a_m[1];
        end else begin
          state <= add_0;
        end
      end

      add_0:
      begin
        z_e <= a_e;
        if (a_s == b_s) begin
          sum <= a_m + b_m;
          z_s <= a_s;
        end else begin
          if (a_m >= b_m) begin
            sum <= a_m - b_m;
            z_s <= a_s;
          end else begin
            sum <= b_m - a_m;
            z_s <= b_s;
          end
        end
        state <= add_1;
      end

      add_1:
      begin
        if (sum[27]) begin
          z_m <= sum[27:4];
          guard <= sum[3];
          round_bit <= sum[2];
          sticky <= sum[1] | sum[0];
          z_e <= z_e + 1;
        end else begin
          z_m <= sum[26:3];
          guard <= sum[2];
          round_bit <= sum[1];
          sticky <= sum[0];
        end
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0 && $signed(z_e) > -126) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        if ($signed(z_e) == -126 && z_m[23:0] == 24'h0) begin
          z[31] <= 1'b0; // FIX SIGN BUG: -a + a = +0.
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule


//IEEE Floating Point Multiplier (Single Precision)
//Copyright (C) Jonathan P Dawson 2013
//2013-12-12
module multiplier_9 (
	input_a,
        input_b,
        input_a_stb,
        input_b_stb,
        output_z_ack,
        clk,
        rst,
        output_z,
        output_z_stb,
        input_a_ack,
        input_b_ack);

  input     clk;
  input     rst;

  input     [31:0] input_a;
  input     input_a_stb;
  output    input_a_ack;

  input     [31:0] input_b;
  input     input_b_stb;
  output    input_b_ack;

  output    [31:0] output_z;
  output    output_z_stb;
  input     output_z_ack;

  reg       s_output_z_stb;
  reg       [31:0] s_output_z;
  reg       s_input_a_ack;
  reg       s_input_b_ack;

  reg       [3:0] state;
  parameter get_a         = 4'd0,
            get_b         = 4'd1,
            unpack        = 4'd2,
            special_cases = 4'd3,
            normalise_a   = 4'd4,
            normalise_b   = 4'd5,
            multiply_0    = 4'd6,
            multiply_1    = 4'd7,
            normalise_1   = 4'd8,
            normalise_2   = 4'd9,
            round         = 4'd10,
            pack          = 4'd11,
            put_z         = 4'd12;

  reg       [31:0] a, b, z;
  reg       [23:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [47:0] product;

  always @(posedge clk)
  begin

    case(state)

      get_a:
      begin
        s_input_a_ack <= 1;
        if (s_input_a_ack && input_a_stb) begin
          a <= input_a;
          s_input_a_ack <= 0;
          state <= get_b;
        end
      end

      get_b:
      begin
        s_input_b_ack <= 1;
        if (s_input_b_ack && input_b_stb) begin
          b <= input_b;
          s_input_b_ack <= 0;
          state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[22 : 0];
        b_m <= b[22 : 0];
        a_e <= a[30 : 23] - 127;
        b_e <= b[30 : 23] - 127;
        a_s <= a[31];
        b_s <= b[31];
        state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[31] <= 1;
          z[30:23] <= 255;
          z[22] <= 1;
          z[21:0] <= 0;
          state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 255;
          z[22:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[31] <= 1;
            z[30:23] <= 255;
            z[22] <= 1;
            z[21:0] <= 0;
          end
          state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[31] <= a_s ^ b_s;
          z[30:23] <= 0;
          z[22:0] <= 0;
          state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[23] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[23] <= 1;
          end
          state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[23]) begin
          state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[23]) begin
          state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m;
        state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[47:24];
        guard <= product[23];
        round_bit <= product[22];
        sticky <= (product[21:0] != 0);
        state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[23] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 24'hffffff) begin
            z_e <=z_e + 1;
          end
        end
        state <= pack;
      end

      pack:
      begin
        z[22 : 0] <= z_m[22:0];
        z[30 : 23] <= z_e[7:0] + 127;
        z[31] <= z_s;
        if ($signed(z_e) == -126 && z_m[23] == 0) begin
          z[30 : 23] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[22 : 0] <= 0;
          z[30 : 23] <= 255;
          z[31] <= z_s;
        end
        state <= put_z;
      end

      put_z:
      begin
        s_output_z_stb <= 1;
        s_output_z <= z;
        if (s_output_z_stb && output_z_ack) begin
          s_output_z_stb <= 0;
          state <= get_a;
        end
      end

    endcase

    if (rst == 1) begin
      state <= get_a;
      s_input_a_ack <= 0;
      s_input_b_ack <= 0;
      s_output_z_stb <= 0;
    end

  end
  assign input_a_ack = s_input_a_ack;
  assign input_b_ack = s_input_b_ack;
  assign output_z_stb = s_output_z_stb;
  assign output_z = s_output_z;
endmodule

